-- cordic_inst0.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cordic_inst0 is
	port (
		a      : in  std_logic_vector(12 downto 0) := (others => '0'); --      a.a
		areset : in  std_logic                     := '0';             -- areset.reset
		c      : out std_logic_vector(9 downto 0);                     --      c.c
		clk    : in  std_logic                     := '0';             --    clk.clk
		s      : out std_logic_vector(9 downto 0)                      --      s.s
	);
end entity cordic_inst0;

architecture rtl of cordic_inst0 is
	component cordic_inst0_CORDIC_0 is
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			areset : in  std_logic                     := 'X';             -- reset
			a      : in  std_logic_vector(12 downto 0) := (others => 'X'); -- a
			c      : out std_logic_vector(9 downto 0);                     -- c
			s      : out std_logic_vector(9 downto 0)                      -- s
		);
	end component cordic_inst0_CORDIC_0;

begin

	cordic_0 : component cordic_inst0_CORDIC_0
		port map (
			clk    => clk,    --    clk.clk
			areset => areset, -- areset.reset
			a      => a,      --      a.a
			c      => c,      --      c.c
			s      => s       --      s.s
		);

end architecture rtl; -- of cordic_inst0
