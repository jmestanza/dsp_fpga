// unnamed.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module unnamed (
		input  wire [12:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [9:0]  c,      //      c.c
		input  wire        clk,    //    clk.clk
		output wire [9:0]  s       //      s.s
	);

	unnamed_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
