// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
// CREATED		"Thu Nov 26 13:10:01 2020"

module PWMyLED(
	Clock,
	cout
);


input wire	Clock;
output wire	cout;

wire	[19:0] qout;
wire	SYNTHESIZED_WIRE_0;





pwm_ip	b2v_inst(
	.inclk0(Clock),
	.c0(SYNTHESIZED_WIRE_0));


upcounter20b	b2v_inst1(
	.clock(SYNTHESIZED_WIRE_0),
	.q(qout));

assign	cout = qout[19];

endmodule
