-- unnamed.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unnamed is
	port (
		a      : in  std_logic_vector(12 downto 0) := (others => '0'); --      a.a
		areset : in  std_logic                     := '0';             -- areset.reset
		c      : out std_logic_vector(9 downto 0);                     --      c.c
		clk    : in  std_logic                     := '0';             --    clk.clk
		s      : out std_logic_vector(9 downto 0)                      --      s.s
	);
end entity unnamed;

architecture rtl of unnamed is
	component unnamed_CORDIC_0 is
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			areset : in  std_logic                     := 'X';             -- reset
			a      : in  std_logic_vector(12 downto 0) := (others => 'X'); -- a
			c      : out std_logic_vector(9 downto 0);                     -- c
			s      : out std_logic_vector(9 downto 0)                      -- s
		);
	end component unnamed_CORDIC_0;

begin

	cordic_0 : component unnamed_CORDIC_0
		port map (
			clk    => clk,    --    clk.clk
			areset => areset, -- areset.reset
			a      => a,      --      a.a
			c      => c,      --      c.c
			s      => s       --      s.s
		);

end architecture rtl; -- of unnamed
