module sonic_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [107:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		12'b000000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b000000001110: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111100010011111;
		12'b000000001111: color_data = 108'b111111111111111111111111111111111111111111111111100010011111111111111111111111111111111011101111011110001111;
		12'b000000010000: color_data = 108'b111111111111111111111111111111111111111111111111011110001111111111111111111111111111100010011111011110001111;
		12'b000000010001: color_data = 108'b111111111111111111111111111111111111111111111111011110001111111111111111111111111111011110001111011110001111;
		12'b000000010010: color_data = 108'b111111111111111111111111111111111111111111111111011110001111111111111111111111111111011110001111011110001111;
		12'b000000010011: color_data = 108'b111111111111111111111111111111111111111111111111011110001111111111111111111111111111011110001111011110001111;
		12'b000000010100: color_data = 108'b111111111111111111111111111111111111111111111111011110001111111111111111111111111111011110001111100110101111;
		12'b000000010101: color_data = 108'b111111111111111111111111111111111111111111111111100110101111111111111111111111111111011110001111111111111111;
		12'b000000010110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110101111111111111111;
		12'b000000010111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000011111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001111;
		12'b000001001000: color_data = 108'b111111111111111111111111111111111111111111111111110011001111111111111111111111111111111111111111101110111111;
		12'b000001001001: color_data = 108'b111111111111111111111111111111111111111111111111101110111111111111111111111111111111110011001111101110111111;
		12'b000001001010: color_data = 108'b111111111111111111111111111111111111111111111111101110111111111111111111111111111111101110111111101110111111;
		12'b000001001011: color_data = 108'b111111111111111111111111111111111111111111111111101110111111111111111111111111111111101110111111101110111111;
		12'b000001001100: color_data = 108'b111111111111111111111111111111111111111111111111101110111111111111111111111111111111101110111111101111001111;
		12'b000001001101: color_data = 108'b111111111111111111111111111011101111111111111111101111001111111111111111111111111111101110111111101010111111;
		12'b000001001110: color_data = 108'b111011101111111111111111100010011111111111111111101010111111111111111111111111111111101111001111001101011111;
		12'b000001001111: color_data = 108'b100010011111111011101111011110001111111111111111001101011111111111111111111111111111101010111111001001001111;
		12'b000001010000: color_data = 108'b011110001111100010011111011110001111111111111111001001001111111111111111111111111111001101011111001001001111;
		12'b000001010001: color_data = 108'b011110001111011110001111011110001111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000001010010: color_data = 108'b011110001111011110001111011110001111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000001010011: color_data = 108'b011110001111011110001111011110001111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000001010100: color_data = 108'b011110001111011110001111100110101111111111111111001001001111111111111111111111111111001001001111010001101111;
		12'b000001010101: color_data = 108'b100110101111011110001111111111111111111111111111010001101111111111111111111111111111001001001111101110111111;
		12'b000001010110: color_data = 108'b111111111111100110101111111111111111111111111111101110111111111111111111111111111111010001101111101110111111;
		12'b000001010111: color_data = 108'b111111111111111111111111111111111111111111111111101110111111111111111111111111111111101110111111101110111111;
		12'b000001011000: color_data = 108'b111111111111111111111111111111111111111111111111101110111111111111111111111111111111101110111111110011001111;
		12'b000001011001: color_data = 108'b111111111111111111111111111111111111111111111111110011001111111111111111111111111111101110111111111011111111;
		12'b000001011010: color_data = 108'b111111111111111111111111111111111111111111111111111011111111111111111111111111111111110011001111111111111111;
		12'b000001011011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111;
		12'b000001011100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001011101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001011110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001011111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110;
		12'b000010000101: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111111011101110;
		12'b000010000110: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111011101110110111011110;
		12'b000010000111: color_data = 108'b111111111111111111111111110011001111111111111111110111011110111111111111111111111111111011101110010101101111;
		12'b000010001000: color_data = 108'b110011001111111111111111101110111111111111111111010101101111111111111111111111111111110111011110001001001111;
		12'b000010001001: color_data = 108'b101110111111110011001111101110111111111111111111001001001111111111111111111111111111010101101111001001001111;
		12'b000010001010: color_data = 108'b101110111111101110111111101110111111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000010001011: color_data = 108'b101110111111101110111111101110111111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000010001100: color_data = 108'b101110111111101110111111101111001111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000010001101: color_data = 108'b101111001111101110111111101010111111111111111111001001001111111111111111111011101111001001001111001001001111;
		12'b000010001110: color_data = 108'b101010111111101111001111001101011111111011101111001001001111111111111111100010011111001001001111001001001111;
		12'b000010001111: color_data = 108'b001101011111101010111111001001001111100010011111001001001111111011101111011110001111001001001111001001001111;
		12'b000010010000: color_data = 108'b001001001111001101011111001001001111011110001111001001001111100010011111011110001111001001001111001001001111;
		12'b000010010001: color_data = 108'b001001001111001001001111001001001111011110001111001001001111011110001111011110001111001001001111001001001111;
		12'b000010010010: color_data = 108'b001001001111001001001111001001001111011110001111001001001111011110001111011110001111001001001111001101011111;
		12'b000010010011: color_data = 108'b001001001111001001001111001001001111011110001111001101011111011110001111011110001111001001001111001101011111;
		12'b000010010100: color_data = 108'b001001001111001001001111010001101111011110001111001101011111011110001111100110101111001101011111001101011111;
		12'b000010010101: color_data = 108'b010001101111001001001111101110111111100110101111001101011111011110001111111111111111001101011111001001001111;
		12'b000010010110: color_data = 108'b101110111111010001101111101110111111111111111111001001001111100110101111111111111111001101011111001001001111;
		12'b000010010111: color_data = 108'b101110111111101110111111101110111111111111111111001001001111111111111111111111111111001001001111001001001111;
		12'b000010011000: color_data = 108'b101110111111101110111111110011001111111111111111001001001111111111111111111111111111001001001111010101101111;
		12'b000010011001: color_data = 108'b110011001111101110111111111011111111111111111111010101101111111111111111111111111111001001001111110111011111;
		12'b000010011010: color_data = 108'b111011111111110011001111111111111111111111111111110111011111111111111111111111111111010101101111111011101111;
		12'b000010011011: color_data = 108'b111111111111111011111111111111111111111111111111111011101111111111111111111111111111110111011111111011101111;
		12'b000010011100: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111011101111111111111111;
		12'b000010011101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111;
		12'b000010011110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010011111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110;
		12'b000010100010: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111111011101110;
		12'b000010100011: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111011101110111111111111;
		12'b000010100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111;
		12'b000010100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011000100: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111111111111111111111111100110011100;
		12'b000011000101: color_data = 108'b111011101110111111111111111011101110111111111111100110011100111111111111111111111111111111111111001101001010;
		12'b000011000110: color_data = 108'b111011101110111011101110110111011110111111111111001101001010111111111111111111111111100110011100001101001010;
		12'b000011000111: color_data = 108'b110111011110111011101110010101101111111111111111001101001010111111111111110011001111001101001010001000111010;
		12'b000011001000: color_data = 108'b010101101111110111011110001001001111110011001111001000111010111111111111101110111111001101001010000100101010;
		12'b000011001001: color_data = 108'b001001001111010101101111001001001111101110111111000100101010110011001111101110111111001000111010000100111011;
		12'b000011001010: color_data = 108'b001001001111001001001111001001001111101110111111000100111011101110111111101110111111000100101010001001001111;
		12'b000011001011: color_data = 108'b001001001111001001001111001001001111101110111111001001001111101110111111101110111111000100111011001001001111;
		12'b000011001100: color_data = 108'b001001001111001001001111001001001111101110111111001001001111101110111111101111001111001001001111001001001111;
		12'b000011001101: color_data = 108'b001001001111001001001111001001001111101111001111001001001111101110111111101010111111001001001111001001001111;
		12'b000011001110: color_data = 108'b001001001111001001001111001001001111101010111111001001001111101111001111001101011111001001001111001001001111;
		12'b000011001111: color_data = 108'b001001001111001001001111001001001111001101011111001001001111101010111111001001001111001001001111001001001111;
		12'b000011010000: color_data = 108'b001001001111001001001111001001001111001001001111001001001111001101011111001001001111001001001111001001001111;
		12'b000011010001: color_data = 108'b001001001111001001001111001001001111001001001111001001001111001001001111001001001111001001001111001001001111;
		12'b000011010010: color_data = 108'b001001001111001001001111001101011111001001001111001001001111001001001111001001001111001001001111000100111011;
		12'b000011010011: color_data = 108'b001101011111001001001111001101011111001001001111000100111011001001001111001001001111001001001111000100111010;
		12'b000011010100: color_data = 108'b001101011111001101011111001101011111001001001111000100111010001001001111010001101111000100111011001000111011;
		12'b000011010101: color_data = 108'b001101011111001101011111001001001111010001101111001000111011001001001111101110111111000100111010001101011111;
		12'b000011010110: color_data = 108'b001001001111001101011111001001001111101110111111001101011111010001101111101110111111001000111011001101011111;
		12'b000011010111: color_data = 108'b001001001111001001001111001001001111101110111111001101011111101110111111101110111111001101011111001101011111;
		12'b000011011000: color_data = 108'b001001001111001001001111010101101111101110111111001101011111101110111111110011001111001101011111001101011111;
		12'b000011011001: color_data = 108'b010101101111001001001111110111011111110011001111001101011111101110111111111011111111001101011111010001101111;
		12'b000011011010: color_data = 108'b110111011111010101101111111011101111111011111111010001101111110011001111111111111111001101011111010001101111;
		12'b000011011011: color_data = 108'b111011101111110111011111111011101111111111111111010001101111111011111111111111111111010001101111100010011111;
		12'b000011011100: color_data = 108'b111011101111111011101111111111111111111111111111100010011111111111111111111111111111010001101111111111111111;
		12'b000011011101: color_data = 108'b111111111111111011101111111111111111111111111111111111111111111111111111111111111111100010011111111111111111;
		12'b000011011110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011011111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110;
		12'b000011100001: color_data = 108'b111111111111111111111111111011101110111111111111111011101110111111111111111111111111111111111111010101101011;
		12'b000011100010: color_data = 108'b111011101110111111111111111011101110111111111111010101101011111111111111111111111111111011101110100110101100;
		12'b000011100011: color_data = 108'b111011101110111011101110111111111111111111111111100110101100111111111111111111111111010101101011111111111111;
		12'b000011100100: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111111111111111111111111100110101100111111111111;
		12'b000011100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100000100: color_data = 108'b111111111111111111111111100110011100111111111111111111111111111111111111111011101110111111111111101110111101;
		12'b000100000101: color_data = 108'b100110011100111111111111001101001010111011101110101110111101111111111111111011101110111111111111100010011100;
		12'b000100000110: color_data = 108'b001101001010100110011100001101001010111011101110100010011100111011101110110111011110101110111101100010011100;
		12'b000100000111: color_data = 108'b001101001010001101001010001000111010110111011110100010011100111011101110010101101111100010011100100010011100;
		12'b000100001000: color_data = 108'b001000111010001101001010000100101010010101101111100010011100110111011110001001001111100010011100010101101010;
		12'b000100001001: color_data = 108'b000100101010001000111010000100111011001001001111010101101010010101101111001001001111100010011100000100101001;
		12'b000100001010: color_data = 108'b000100111011000100101010001001001111001001001111000100101001001001001111001001001111010101101010000100111011;
		12'b000100001011: color_data = 108'b001001001111000100111011001001001111001001001111000100111011001001001111001001001111000100101001000100111100;
		12'b000100001100: color_data = 108'b001001001111001001001111001001001111001001001111000100111100001001001111001001001111000100111011000100111100;
		12'b000100001101: color_data = 108'b001001001111001001001111001001001111001001001111000100111100001001001111001001001111000100111100001000111100;
		12'b000100001110: color_data = 108'b001001001111001001001111001001001111001001001111001000111100001001001111001001001111000100111100001000111100;
		12'b000100001111: color_data = 108'b001001001111001001001111001001001111001001001111001000111100001001001111001001001111001000111100001001001110;
		12'b000100010000: color_data = 108'b001001001111001001001111001001001111001001001111001001001110001001001111001001001111001000111100001001001111;
		12'b000100010001: color_data = 108'b001001001111001001001111001001001111001001001111001001001111001001001111001001001111001001001110001001001111;
		12'b000100010010: color_data = 108'b001001001111001001001111000100111011001001001111001001001111001001001111001101011111001001001111000100101010;
		12'b000100010011: color_data = 108'b000100111011001001001111000100111010001101011111000100101010001001001111001101011111001001001111010101011001;
		12'b000100010100: color_data = 108'b000100111010000100111011001000111011001101011111010101011001001101011111001101011111000100101010011101101010;
		12'b000100010101: color_data = 108'b001000111011000100111010001101011111001101011111011101101010001101011111001001001111010101011001001001001100;
		12'b000100010110: color_data = 108'b001101011111001000111011001101011111001001001111001001001100001101011111001001001111011101101010001101011111;
		12'b000100010111: color_data = 108'b001101011111001101011111001101011111001001001111001101011111001001001111001001001111001001001100001101101111;
		12'b000100011000: color_data = 108'b001101011111001101011111001101011111001001001111001101101111001001001111010101101111001101011111001101101111;
		12'b000100011001: color_data = 108'b001101011111001101011111010001101111010101101111001101101111001001001111110111011111001101101111001001011111;
		12'b000100011010: color_data = 108'b010001101111001101011111010001101111110111011111001001011111010101101111111011101111001101101111001001011111;
		12'b000100011011: color_data = 108'b010001101111010001101111100010011111111011101111001001011111110111011111111011101111001001011111010101101111;
		12'b000100011100: color_data = 108'b100010011111010001101111111111111111111011101111010101101111111011101111111111111111001001011111100010011111;
		12'b000100011101: color_data = 108'b111111111111100010011111111111111111111111111111100010011111111011101111111111111111010101101111100010011111;
		12'b000100011110: color_data = 108'b111111111111111111111111111111111111111111111111100010011111111111111111111111111111100010011111110011011111;
		12'b000100011111: color_data = 108'b111111111111111111111111111111111111111111111111110011011111111111111111111111111111100010011111110111011110;
		12'b000100100000: color_data = 108'b111111111111111111111111111011101110111111111111110111011110111111111111111111111111110011011111011110001011;
		12'b000100100001: color_data = 108'b111011101110111111111111010101101011111111111111011110001011111111111111111011101110110111011110001000111001;
		12'b000100100010: color_data = 108'b010101101011111011101110100110101100111011101110001000111001111111111111111011101110011110001011100010011100;
		12'b000100100011: color_data = 108'b100110101100010101101011111111111111111011101110100010011100111011101110111111111111001000111001111111111111;
		12'b000100100100: color_data = 108'b111111111111100110101100111111111111111111111111111111111111111011101110111111111111100010011100111111111111;
		12'b000100100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101000100: color_data = 108'b111111111111111111111111101110111101111111111111111111111111111111111111100110011100111111111111111111111111;
		12'b000101000101: color_data = 108'b101110111101111111111111100010011100100110011100111111111111111111111111001101001010111111111111111111111111;
		12'b000101000110: color_data = 108'b100010011100101110111101100010011100001101001010111111111111100110011100001101001010111111111111111111111111;
		12'b000101000111: color_data = 108'b100010011100100010011100100010011100001101001010111111111111001101001010001000111010111111111111111111111111;
		12'b000101001000: color_data = 108'b100010011100100010011100010101101010001000111010111111111111001101001010000100101010111111111111101010101101;
		12'b000101001001: color_data = 108'b010101101010100010011100000100101001000100101010101010101101001000111010000100111011111111111111010001011010;
		12'b000101001010: color_data = 108'b000100101001010101101010000100111011000100111011010001011010000100101010001001001111101010101101010001011010;
		12'b000101001011: color_data = 108'b000100111011000100101001000100111100001001001111010001011010000100111011001001001111010001011010010001011010;
		12'b000101001100: color_data = 108'b000100111100000100111011000100111100001001001111010001011010001001001111001001001111010001011010001101001001;
		12'b000101001101: color_data = 108'b000100111100000100111100001000111100001001001111001101001001001001001111001001001111010001011010000100101000;
		12'b000101001110: color_data = 108'b001000111100000100111100001000111100001001001111000100101000001001001111001001001111001101001001000100101000;
		12'b000101001111: color_data = 108'b001000111100001000111100001001001110001001001111000100101000001001001111001001001111000100101000001000111100;
		12'b000101010000: color_data = 108'b001001001110001000111100001001001111001001001111001000111100001001001111001001001111000100101000001000111110;
		12'b000101010001: color_data = 108'b001001001111001001001110001001001111001001001111001000111110001001001111001001001111001000111100001000111101;
		12'b000101010010: color_data = 108'b001001001111001001001111000100101010001001001111001000111101001001001111000100111011001000111110001100111001;
		12'b000101010011: color_data = 108'b000100101010001001001111010101011001000100111011001100111001001001001111000100111010001000111101101010001001;
		12'b000101010100: color_data = 108'b010101011001000100101010011101101010000100111010101010001001000100111011001000111011001100111001110110101001;
		12'b000101010101: color_data = 108'b011101101010010101011001001001001100001000111011110110101001000100111010001101011111101010001001010101011001;
		12'b000101010110: color_data = 108'b001001001100011101101010001101011111001101011111010101011001001000111011001101011111110110101001001101011100;
		12'b000101010111: color_data = 108'b001101011111001001001100001101101111001101011111001101011100001101011111001101011111010101011001001101011111;
		12'b000101011000: color_data = 108'b001101101111001101011111001101101111001101011111001101011111001101011111001101011111001101011100001101101111;
		12'b000101011001: color_data = 108'b001101101111001101101111001001011111001101011111001101101111001101011111010001101111001101011111010001101111;
		12'b000101011010: color_data = 108'b001001011111001101101111001001011111010001101111010001101111001101011111010001101111001101101111001101101111;
		12'b000101011011: color_data = 108'b001001011111001001011111010101101111010001101111001101101111010001101111100010011111010001101111001101011111;
		12'b000101011100: color_data = 108'b010101101111001001011111100010011111100010011111001101011111010001101111111111111111001101101111001001001111;
		12'b000101011101: color_data = 108'b100010011111010101101111100010011111111111111111001001001111100010011111111111111111001101011111001001001111;
		12'b000101011110: color_data = 108'b100010011111100010011111110011011111111111111111001001001111111111111111111111111111001001001111100010011111;
		12'b000101011111: color_data = 108'b110011011111100010011111110111011110111111111111100010011111111111111111111111111111001001001111100110011101;
		12'b000101100000: color_data = 108'b110111011110110011011111011110001011111111111111100110011101111111111111111011101110100010011111000100101001;
		12'b000101100001: color_data = 108'b011110001011110111011110001000111001111011101110000100101001111111111111010101101011100110011101000100101001;
		12'b000101100010: color_data = 108'b001000111001011110001011100010011100010101101011000100101001111011101110100110101100000100101001100010011100;
		12'b000101100011: color_data = 108'b100010011100001000111001111111111111100110101100100010011100010101101011111111111111000100101001111111111111;
		12'b000101100100: color_data = 108'b111111111111100010011100111111111111111111111111111111111111100110101100111111111111100010011100111111111111;
		12'b000101100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111101110111101111111111111111111111111;
		12'b000110000101: color_data = 108'b111111111111111111111111111111111111101110111101111111111111111111111111100010011100111111111111111111111111;
		12'b000110000110: color_data = 108'b111111111111111111111111111111111111100010011100111111111111101110111101100010011100111111111111111111111111;
		12'b000110000111: color_data = 108'b111111111111111111111111111111111111100010011100111111111111100010011100100010011100111111111111111111111111;
		12'b000110001000: color_data = 108'b111111111111111111111111101010101101100010011100111111111111100010011100010101101010111111111111111011101111;
		12'b000110001001: color_data = 108'b101010101101111111111111010001011010010101101010111011101111100010011100000100101001111111111111111011101110;
		12'b000110001010: color_data = 108'b010001011010101010101101010001011010000100101001111011101110010101101010000100111011111011101111111011101110;
		12'b000110001011: color_data = 108'b010001011010010001011010010001011010000100111011111011101110000100101001000100111100111011101110111011101111;
		12'b000110001100: color_data = 108'b010001011010010001011010001101001001000100111100111011101111000100111011000100111100111011101110100110101100;
		12'b000110001101: color_data = 108'b001101001001010001011010000100101000000100111100100110101100000100111100001000111100111011101111000100101001;
		12'b000110001110: color_data = 108'b000100101000001101001001000100101000001000111100000100101001000100111100001000111100100110101100000100101001;
		12'b000110001111: color_data = 108'b000100101000000100101000001000111100001000111100000100101001001000111100001001001110000100101001000100101001;
		12'b000110010000: color_data = 108'b001000111100000100101000001000111110001001001110000100101001001000111100001001001111000100101001000100101001;
		12'b000110010001: color_data = 108'b001000111110001000111100001000111101001001001111000100101001001001001110001001001111000100101001001000101001;
		12'b000110010010: color_data = 108'b001000111101001000111110001100111001001001001111001000101001001001001111000100101010000100101001100101100110;
		12'b000110010011: color_data = 108'b001100111001001000111101101010001001000100101010100101100110001001001111010101011001001000101001110110100111;
		12'b000110010100: color_data = 108'b101010001001001100111001110110101001010101011001110110100111000100101010011101101010100101100110111111001010;
		12'b000110010101: color_data = 108'b110110101001101010001001010101011001011101101010111111001010010101011001001001001100110110100111111010111010;
		12'b000110010110: color_data = 108'b010101011001110110101001001101011100001001001100111010111010011101101010001101011111111111001010010101011001;
		12'b000110010111: color_data = 108'b001101011100010101011001001101011111001101011111010101011001001001001100001101101111111010111010001001001100;
		12'b000110011000: color_data = 108'b001101011111001101011100001101101111001101101111001001001100001101011111001101101111010101011001001101101111;
		12'b000110011001: color_data = 108'b001101101111001101011111010001101111001101101111001101101111001101101111001001011111001001001100010101111111;
		12'b000110011010: color_data = 108'b010001101111001101101111001101101111001001011111010101111111001101101111001001011111001101101111010001101111;
		12'b000110011011: color_data = 108'b001101101111010001101111001101011111001001011111010001101111001001011111010101101111010101111111001101101111;
		12'b000110011100: color_data = 108'b001101011111001101101111001001001111010101101111001101101111001001011111100010011111010001101111001101101111;
		12'b000110011101: color_data = 108'b001001001111001101011111001001001111100010011111001101101111010101101111100010011111001101101111001101101111;
		12'b000110011110: color_data = 108'b001001001111001001001111100010011111100010011111001101101111100010011111110011011111001101101111001101011111;
		12'b000110011111: color_data = 108'b100010011111001001001111100110011101110011011111001101011111100010011111110111011110001101101111001001001101;
		12'b000110100000: color_data = 108'b100110011101100010011111000100101001110111011110001001001101110011011111011110001011001101011111000100101001;
		12'b000110100001: color_data = 108'b000100101001100110011101000100101001011110001011000100101001110111011110001000111001001001001101000100101001;
		12'b000110100010: color_data = 108'b000100101001000100101001100010011100001000111001000100101001011110001011100010011100000100101001100010011100;
		12'b000110100011: color_data = 108'b100010011100000100101001111111111111100010011100100010011100001000111001111111111111000100101001111111111111;
		12'b000110100100: color_data = 108'b111111111111100010011100111111111111111111111111111111111111100010011100111111111111100010011100111111111111;
		12'b000110100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b000111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111001000: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111101010101101111111111111111111111111;
		12'b000111001001: color_data = 108'b111011101111111111111111111011101110101010101101111111111111111111111111010001011010111111111111111111111111;
		12'b000111001010: color_data = 108'b111011101110111011101111111011101110010001011010111111111111101010101101010001011010111111111111111111111111;
		12'b000111001011: color_data = 108'b111011101110111011101110111011101111010001011010111111111111010001011010010001011010111111111111111111111111;
		12'b000111001100: color_data = 108'b111011101111111011101110100110101100010001011010111111111111010001011010001101001001111111111111111011101110;
		12'b000111001101: color_data = 108'b100110101100111011101111000100101001001101001001111011101110010001011010000100101000111111111111101010111101;
		12'b000111001110: color_data = 108'b000100101001100110101100000100101001000100101000101010111101001101001001000100101000111011101110001000111001;
		12'b000111001111: color_data = 108'b000100101001000100101001000100101001000100101000001000111001000100101000001000111100101010111101000100111100;
		12'b000111010000: color_data = 108'b000100101001000100101001000100101001001000111100000100111100000100101000001000111110001000111001001000111100;
		12'b000111010001: color_data = 108'b000100101001000100101001001000101001001000111110001000111100001000111100001000111101000100111100001000101000;
		12'b000111010010: color_data = 108'b001000101001000100101001100101100110001000111101001000101000001000111110001100111001001000111100100101100101;
		12'b000111010011: color_data = 108'b100101100110001000101001110110100111001100111001100101100101001000111101101010001001001000101000111010100111;
		12'b000111010100: color_data = 108'b110110100111100101100110111111001010101010001001111010100111001100111001110110101001100101100101111111001010;
		12'b000111010101: color_data = 108'b111111001010110110100111111010111010110110101001111111001010101010001001010101011001111010100111111111001001;
		12'b000111010110: color_data = 108'b111010111010111111001010010101011001010101011001111111001001110110101001001101011100111111001010110110101001;
		12'b000111010111: color_data = 108'b010101011001111010111010001001001100001101011100110110101001010101011001001101011111111111001001100001111100;
		12'b000111011000: color_data = 108'b001001001100010101011001001101101111001101011111100001111100001101011100001101101111110110101001001101011111;
		12'b000111011001: color_data = 108'b001101101111001001001100010101111111001101101111001101011111001101011111010001101111100001111100010101111111;
		12'b000111011010: color_data = 108'b010101111111001101101111010001101111010001101111010101111111001101101111001101101111001101011111010101111111;
		12'b000111011011: color_data = 108'b010001101111010101111111001101101111001101101111010101111111010001101111001101011111010101111111010101111111;
		12'b000111011100: color_data = 108'b001101101111010001101111001101101111001101011111010101111111001101101111001001001111010101111111010101111111;
		12'b000111011101: color_data = 108'b001101101111001101101111001101101111001001001111010101111111001101011111001001001111010101111111001101101111;
		12'b000111011110: color_data = 108'b001101101111001101101111001101011111001001001111001101101111001001001111100010011111010101111111001101011111;
		12'b000111011111: color_data = 108'b001101011111001101101111001001001101100010011111001101011111001001001111100110011101001101101111001101011111;
		12'b000111100000: color_data = 108'b001001001101001101011111000100101001100110011101001101011111100010011111000100101001001101011111001000111101;
		12'b000111100001: color_data = 108'b000100101001001001001101000100101001000100101001001000111101100110011101000100101001001101011111000100101001;
		12'b000111100010: color_data = 108'b000100101001000100101001100010011100000100101001000100101001000100101001100010011100001000111101100010011100;
		12'b000111100011: color_data = 108'b100010011100000100101001111111111111100010011100100010011100000100101001111111111111000100101001111111111111;
		12'b000111100100: color_data = 108'b111111111111100010011100111111111111111111111111111111111111100010011100111111111111100010011100111111111111;
		12'b000111100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b000111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111;
		12'b001000001001: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111111111111111011101110111111111111111111111111;
		12'b001000001010: color_data = 108'b111111111111111111111111111111111111111011101110111111111111111011101111111011101110111111111111111111111111;
		12'b001000001011: color_data = 108'b111111111111111111111111111111111111111011101110111111111111111011101110111011101111111111111111111111111111;
		12'b001000001100: color_data = 108'b111111111111111111111111111011101110111011101111111111111111111011101110100110101100111111111111110111011111;
		12'b001000001101: color_data = 108'b111011101110111111111111101010111101100110101100110111011111111011101111000100101001111111111111100010011111;
		12'b001000001110: color_data = 108'b101010111101111011101110001000111001000100101001100010011111100110101100000100101001110111011111001001001100;
		12'b001000001111: color_data = 108'b001000111001101010111101000100111100000100101001001001001100000100101001000100101001100010011111001001001110;
		12'b001000010000: color_data = 108'b000100111100001000111001001000111100000100101001001001001110000100101001000100101001001001001100001000111101;
		12'b001000010001: color_data = 108'b001000111100000100111100001000101000000100101001001000111101000100101001001000101001001001001110001000101000;
		12'b001000010010: color_data = 108'b001000101000001000111100100101100101001000101001001000101000000100101001100101100110001000111101100101100101;
		12'b001000010011: color_data = 108'b100101100101001000101000111010100111100101100110100101100101001000101001110110100111001000101000110110010110;
		12'b001000010100: color_data = 108'b111010100111100101100101111111001010110110100111110110010110100101100110111111001010100101100101110110101001;
		12'b001000010101: color_data = 108'b111111001010111010100111111111001001111111001010110110101001110110100111111010111010110110010110101010011100;
		12'b001000010110: color_data = 108'b111111001001111111001010110110101001111010111010101010011100111111001010010101011001110110101001101010011100;
		12'b001000010111: color_data = 108'b110110101001111111001001100001111100010101011001101010011100111010111010001001001100101010011100011101111110;
		12'b001000011000: color_data = 108'b100001111100110110101001001101011111001001001100011101111110010101011001001101101111101010011100010001101111;
		12'b001000011001: color_data = 108'b001101011111100001111100010101111111001101101111010001101111001001001100010101111111011101111110011001111111;
		12'b001000011010: color_data = 108'b010101111111001101011111010101111111010101111111011001111111001101101111010001101111010001101111011001111111;
		12'b001000011011: color_data = 108'b010101111111010101111111010101111111010001101111011001111111010101111111001101101111011001111111011001111111;
		12'b001000011100: color_data = 108'b010101111111010101111111010101111111001101101111011001111111010001101111001101101111011001111111011001111111;
		12'b001000011101: color_data = 108'b010101111111010101111111001101101111001101101111011001111111001101101111001101101111011001111111010001111111;
		12'b001000011110: color_data = 108'b001101101111010101111111001101011111001101101111010001111111001101101111001101011111011001111111001101101111;
		12'b001000011111: color_data = 108'b001101011111001101101111001101011111001101011111001101101111001101101111001001001101010001111111001101011111;
		12'b001000100000: color_data = 108'b001101011111001101011111001000111101001001001101001101011111001101011111000100101001001101101111001001011111;
		12'b001000100001: color_data = 108'b001000111101001101011111000100101001000100101001001001011111001001001101000100101001001101011111001000111100;
		12'b001000100010: color_data = 108'b000100101001001000111101100010011100000100101001001000111100000100101001100010011100001001011111100110011101;
		12'b001000100011: color_data = 108'b100010011100000100101001111111111111100010011100100110011101000100101001111111111111001000111100111111111111;
		12'b001000100100: color_data = 108'b111111111111100010011100111111111111111111111111111111111111100010011100111111111111100110011101111111111111;
		12'b001000100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b001001001010: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111110111011111;
		12'b001001001011: color_data = 108'b111111111111111111111111111111111111111111111111110111011111111111111111111111111111111011101111110111011111;
		12'b001001001100: color_data = 108'b111111111111111111111111110111011111111111111111110111011111111111111111111011101110110111011111100110101111;
		12'b001001001101: color_data = 108'b110111011111111111111111100010011111111011101110100110101111111111111111101010111101110111011111001001001111;
		12'b001001001110: color_data = 108'b100010011111110111011111001001001100101010111101001001001111111011101110001000111001100110101111001001001110;
		12'b001001001111: color_data = 108'b001001001100100010011111001001001110001000111001001001001110101010111101000100111100001001001111001001001111;
		12'b001001010000: color_data = 108'b001001001110001001001100001000111101000100111100001001001111001000111001001000111100001001001110001000111110;
		12'b001001010001: color_data = 108'b001000111101001001001110001000101000001000111100001000111110000100111100001000101000001001001111001000111010;
		12'b001001010010: color_data = 108'b001000101000001000111101100101100101001000101000001000111010001000111100100101100101001000111110100001100111;
		12'b001001010011: color_data = 108'b100101100101001000101000110110010110100101100101100001100111001000101000111010100111001000111010101001110110;
		12'b001001010100: color_data = 108'b110110010110100101100101110110101001111010100111101001110110100101100101111111001010100001100111100001111001;
		12'b001001010101: color_data = 108'b110110101001110110010110101010011100111111001010100001111001111010100111111111001001101001110110001101101111;
		12'b001001010110: color_data = 108'b101010011100110110101001101010011100111111001001001101101111111111001010110110101001100001111001001101101111;
		12'b001001010111: color_data = 108'b101010011100101010011100011101111110110110101001001101101111111111001001100001111100001101101111010001101111;
		12'b001001011000: color_data = 108'b011101111110101010011100010001101111100001111100010001101111110110101001001101011111001101101111010101111111;
		12'b001001011001: color_data = 108'b010001101111011101111110011001111111001101011111010101111111100001111100010101111111010001101111010101111111;
		12'b001001011010: color_data = 108'b011001111111010001101111011001111111010101111111010101111111001101011111010101111111010101111111010101111111;
		12'b001001011011: color_data = 108'b011001111111011001111111011001111111010101111111010101111111010101111111010101111111010101111111010101111111;
		12'b001001011100: color_data = 108'b011001111111011001111111011001111111010101111111010101111111010101111111010101111111010101111111010101111111;
		12'b001001011101: color_data = 108'b011001111111011001111111010001111111010101111111010101111111010101111111001101101111010101111111011001111111;
		12'b001001011110: color_data = 108'b010001111111011001111111001101101111001101101111011001111111010101111111001101011111010101111111010001101111;
		12'b001001011111: color_data = 108'b001101101111010001111111001101011111001101011111010001101111001101101111001101011111011001111111001101101111;
		12'b001001100000: color_data = 108'b001101011111001101101111001001011111001101011111001101101111001101011111001000111101010001101111001101101111;
		12'b001001100001: color_data = 108'b001001011111001101011111001000111100001000111101001101101111001101011111000100101001001101101111001001001111;
		12'b001001100010: color_data = 108'b001000111100001001011111100110011101000100101001001001001111001000111101100010011100001101101111100110101111;
		12'b001001100011: color_data = 108'b100110011101001000111100111111111111100010011100100110101111000100101001111111111111001001001111111111111111;
		12'b001001100100: color_data = 108'b111111111111100110011101111111111111111111111111111111111111100010011100111111111111100110101111111111111111;
		12'b001001100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010001001: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111110111011111;
		12'b001010001010: color_data = 108'b111011101111111111111111110111011111111111111111110111011111111111111111111111111111111111111111010001011111;
		12'b001010001011: color_data = 108'b110111011111111011101111110111011111111111111111010001011111111111111111111111111111110111011111001101011111;
		12'b001010001100: color_data = 108'b110111011111110111011111100110101111111111111111001101011111111111111111110111011111010001011111001101001111;
		12'b001010001101: color_data = 108'b100110101111110111011111001001001111110111011111001101001111111111111111100010011111001101011111001001001111;
		12'b001010001110: color_data = 108'b001001001111100110101111001001001110100010011111001001001111110111011111001001001100001101001111000100101010;
		12'b001010001111: color_data = 108'b001001001110001001001111001001001111001001001100000100101010100010011111001001001110001001001111001000111101;
		12'b001010010000: color_data = 108'b001001001111001001001110001000111110001001001110001000111101001001001100001000111101000100101010001001001111;
		12'b001010010001: color_data = 108'b001000111110001001001111001000111010001000111101001001001111001001001110001000101000001000111101001001001111;
		12'b001010010010: color_data = 108'b001000111010001000111110100001100111001000101000001001001111001000111101100101100101001001001111001101001111;
		12'b001010010011: color_data = 108'b100001100111001000111010101001110110100101100101001101001111001000101000110110010110001001001111001101011111;
		12'b001010010100: color_data = 108'b101001110110100001100111100001111001110110010110001101011111100101100101110110101001001101001111010001101111;
		12'b001010010101: color_data = 108'b100001111001101001110110001101101111110110101001010001101111110110010110101010011100001101011111001101101111;
		12'b001010010110: color_data = 108'b001101101111100001111001001101101111101010011100001101101111110110101001101010011100010001101111010101111111;
		12'b001010010111: color_data = 108'b001101101111001101101111010001101111101010011100010101111111101010011100011101111110001101101111010001111111;
		12'b001010011000: color_data = 108'b010001101111001101101111010101111111011101111110010001111111101010011100010001101111010101111111001101101111;
		12'b001010011001: color_data = 108'b010101111111010001101111010101111111010001101111001101101111011101111110011001111111010001111111001101101111;
		12'b001010011010: color_data = 108'b010101111111010101111111010101111111011001111111001101101111010001101111011001111111001101101111001101101111;
		12'b001010011011: color_data = 108'b010101111111010101111111010101111111011001111111001101101111011001111111011001111111001101101111001101101111;
		12'b001010011100: color_data = 108'b010101111111010101111111010101111111011001111111001101101111011001111111011001111111001101101111010001101111;
		12'b001010011101: color_data = 108'b010101111111010101111111011001111111011001111111010001101111011001111111010001111111001101101111010101111111;
		12'b001010011110: color_data = 108'b011001111111010101111111010001101111010001111111010101111111011001111111001101101111010001101111010001101111;
		12'b001010011111: color_data = 108'b010001101111011001111111001101101111001101101111010001101111010001111111001101011111010101111111001101101111;
		12'b001010100000: color_data = 108'b001101101111010001101111001101101111001101011111001101101111001101101111001001011111010001101111001101101111;
		12'b001010100001: color_data = 108'b001101101111001101101111001001001111001001011111001101101111001101011111001000111100001101101111001001001111;
		12'b001010100010: color_data = 108'b001001001111001101101111100110101111001000111100001001001111001001011111100110011101001101101111100110101111;
		12'b001010100011: color_data = 108'b100110101111001001001111111111111111100110011101100110101111001000111100111111111111001001001111111111111111;
		12'b001010100100: color_data = 108'b111111111111100110101111111111111111111111111111111111111111100110011101111111111111100110101111111111111111;
		12'b001010100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010011111;
		12'b001011001000: color_data = 108'b111111111111111111111111111111111111111111111111100010011111111111111111111111111111111111111111011001111111;
		12'b001011001001: color_data = 108'b111111111111111111111111110111011111111111111111011001111111111111111111111011101111100010011111010101111111;
		12'b001011001010: color_data = 108'b110111011111111111111111010001011111111011101111010101111111111111111111110111011111011001111111001001001111;
		12'b001011001011: color_data = 108'b010001011111110111011111001101011111110111011111001001001111111011101111110111011111010101111111001001001111;
		12'b001011001100: color_data = 108'b001101011111010001011111001101001111110111011111001001001111110111011111100110101111001001001111001000111110;
		12'b001011001101: color_data = 108'b001101001111001101011111001001001111100110101111001000111110110111011111001001001111001001001111000100111010;
		12'b001011001110: color_data = 108'b001001001111001101001111000100101010001001001111000100111010100110101111001001001110001000111110000100101001;
		12'b001011001111: color_data = 108'b000100101010001001001111001000111101001001001110000100101001001001001111001001001111000100111010001000111101;
		12'b001011010000: color_data = 108'b001000111101000100101010001001001111001001001111001000111101001001001110001000111110000100101001001001001111;
		12'b001011010001: color_data = 108'b001001001111001000111101001001001111001000111110001001001111001001001111001000111010001000111101001101011111;
		12'b001011010010: color_data = 108'b001001001111001001001111001101001111001000111010001101011111001000111110100001100111001001001111010001101111;
		12'b001011010011: color_data = 108'b001101001111001001001111001101011111100001100111010001101111001000111010101001110110001101011111010101111111;
		12'b001011010100: color_data = 108'b001101011111001101001111010001101111101001110110010101111111100001100111100001111001010001101111010001111111;
		12'b001011010101: color_data = 108'b010001101111001101011111001101101111100001111001010001111111101001110110001101101111010101111111001101101111;
		12'b001011010110: color_data = 108'b001101101111010001101111010101111111001101101111001101101111100001111001001101101111010001111111010001101111;
		12'b001011010111: color_data = 108'b010101111111001101101111010001111111001101101111010001101111001101101111010001101111001101101111001101101111;
		12'b001011011000: color_data = 108'b010001111111010101111111001101101111010001101111001101101111001101101111010101111111010001101111010001101111;
		12'b001011011001: color_data = 108'b001101101111010001111111001101101111010101111111010001101111010001101111010101111111001101101111100010011110;
		12'b001011011010: color_data = 108'b001101101111001101101111001101101111010101111111100010011110010101111111010101111111010001101111100110011101;
		12'b001011011011: color_data = 108'b001101101111001101101111001101101111010101111111100110011101010101111111010101111111100010011110011110001110;
		12'b001011011100: color_data = 108'b001101101111001101101111010001101111010101111111011110001110010101111111010101111111100110011101010101111111;
		12'b001011011101: color_data = 108'b010001101111001101101111010101111111010101111111010101111111010101111111011001111111011110001110010001101111;
		12'b001011011110: color_data = 108'b010101111111010001101111010001101111011001111111010001101111010101111111010001101111010101111111010101111111;
		12'b001011011111: color_data = 108'b010001101111010101111111001101101111010001101111010101111111011001111111001101101111010001101111010001111111;
		12'b001011100000: color_data = 108'b001101101111010001101111001101101111001101101111010001111111010001101111001101101111010101111111001101101111;
		12'b001011100001: color_data = 108'b001101101111001101101111001001001111001101101111001101101111001101101111001001001111010001111111001101011111;
		12'b001011100010: color_data = 108'b001001001111001101101111100110101111001001001111001101011111001101101111100110101111001101101111010001101111;
		12'b001011100011: color_data = 108'b100110101111001001001111111111111111100110101111010001101111001001001111111111111111001101011111100010011111;
		12'b001011100100: color_data = 108'b111111111111100110101111111111111111111111111111100010011111100110101111111111111111010001101111111011101111;
		12'b001011100101: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111100010011111111111111111;
		12'b001011100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111;
		12'b001011100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b001100000110: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111101010111111;
		12'b001100000111: color_data = 108'b111111111111111111111111100010011111111111111111101010111111111111111111111111111111111011101111010001011111;
		12'b001100001000: color_data = 108'b100010011111111111111111011001111111111111111111010001011111111111111111111111111111101010111111001001001111;
		12'b001100001001: color_data = 108'b011001111111100010011111010101111111111111111111001001001111111111111111110111011111010001011111001001001111;
		12'b001100001010: color_data = 108'b010101111111011001111111001001001111110111011111001001001111111111111111010001011111001001001111001001001111;
		12'b001100001011: color_data = 108'b001001001111010101111111001001001111010001011111001001001111110111011111001101011111001001001111001001001111;
		12'b001100001100: color_data = 108'b001001001111001001001111001000111110001101011111001001001111010001011111001101001111001001001111001000111101;
		12'b001100001101: color_data = 108'b001000111110001001001111000100111010001101001111001000111101001101011111001001001111001001001111000100101001;
		12'b001100001110: color_data = 108'b000100111010001000111110000100101001001001001111000100101001001101001111000100101010001000111101000100101001;
		12'b001100001111: color_data = 108'b000100101001000100111010001000111101000100101010000100101001001001001111001000111101000100101001001000111101;
		12'b001100010000: color_data = 108'b001000111101000100101001001001001111001000111101001000111101000100101010001001001111000100101001001101011111;
		12'b001100010001: color_data = 108'b001001001111001000111101001101011111001001001111001101011111001000111101001001001111001000111101010001111111;
		12'b001100010010: color_data = 108'b001101011111001001001111010001101111001001001111010001111111001001001111001101001111001101011111100010101111;
		12'b001100010011: color_data = 108'b010001101111001101011111010101111111001101001111100010101111001001001111001101011111010001111111011110011111;
		12'b001100010100: color_data = 108'b010101111111010001101111010001111111001101011111011110011111001101001111010001101111100010101111010101111111;
		12'b001100010101: color_data = 108'b010001111111010101111111001101101111010001101111010101111111001101011111001101101111011110011111001101101111;
		12'b001100010110: color_data = 108'b001101101111010001111111010001101111001101101111001101101111010001101111010101111111010101111111001101101111;
		12'b001100010111: color_data = 108'b010001101111001101101111001101101111010101111111001101101111001101101111010001111111001101101111010001111111;
		12'b001100011000: color_data = 108'b001101101111010001101111010001101111010001111111010001111111010101111111001101101111001101101111011110001110;
		12'b001100011001: color_data = 108'b010001101111001101101111100010011110001101101111011110001110010001111111001101101111010001111111110011001110;
		12'b001100011010: color_data = 108'b100010011110010001101111100110011101001101101111110011001110001101101111001101101111011110001110110111011110;
		12'b001100011011: color_data = 108'b100110011101100010011110011110001110001101101111110111011110001101101111001101101111110011001110101110111110;
		12'b001100011100: color_data = 108'b011110001110100110011101010101111111001101101111101110111110001101101111010001101111110111011110011110001111;
		12'b001100011101: color_data = 108'b010101111111011110001110010001101111010001101111011110001111001101101111010101111111101110111110010001111111;
		12'b001100011110: color_data = 108'b010001101111010101111111010101111111010101111111010001111111010001101111010001101111011110001111010001111111;
		12'b001100011111: color_data = 108'b010101111111010001101111010001111111010001101111010001111111010101111111001101101111010001111111010001101111;
		12'b001100100000: color_data = 108'b010001111111010101111111001101101111001101101111010001101111010001101111001101101111010001111111001101101111;
		12'b001100100001: color_data = 108'b001101101111010001111111001101011111001101101111001101101111001101101111001001001111010001101111001101101111;
		12'b001100100010: color_data = 108'b001101011111001101101111010001101111001001001111001101101111001101101111100110101111001101101111001101011111;
		12'b001100100011: color_data = 108'b010001101111001101011111100010011111100110101111001101011111001001001111111111111111001101101111011001111111;
		12'b001100100100: color_data = 108'b100010011111010001101111111011101111111111111111011001111111100110101111111111111111001101011111111011101111;
		12'b001100100101: color_data = 108'b111011101111100010011111111111111111111111111111111011101111111111111111111111111111011001111111111111111111;
		12'b001100100110: color_data = 108'b111111111111111011101111111111111111111111111111111111111111111111111111111111111111111011101111111111111111;
		12'b001100100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b001101000101: color_data = 108'b111111111111111111111111111011101111111111111111111011101111111111111111111111111111111111111111101110111111;
		12'b001101000110: color_data = 108'b111011101111111111111111101010111111111111111111101110111111111111111111111111111111111011101111001101001111;
		12'b001101000111: color_data = 108'b101010111111111011101111010001011111111111111111001101001111111111111111100010011111101110111111001001001111;
		12'b001101001000: color_data = 108'b010001011111101010111111001001001111100010011111001001001111111111111111011001111111001101001111001001001111;
		12'b001101001001: color_data = 108'b001001001111010001011111001001001111011001111111001001001111100010011111010101111111001001001111001001001111;
		12'b001101001010: color_data = 108'b001001001111001001001111001001001111010101111111001001001111011001111111001001001111001001001111001001001111;
		12'b001101001011: color_data = 108'b001001001111001001001111001001001111001001001111001001001111010101111111001001001111001001001111001001001111;
		12'b001101001100: color_data = 108'b001001001111001001001111001000111101001001001111001001001111001001001111001000111110001001001111001000111101;
		12'b001101001101: color_data = 108'b001000111101001001001111000100101001001000111110001000111101001001001111000100111010001001001111000100101001;
		12'b001101001110: color_data = 108'b000100101001001000111101000100101001000100111010000100101001001000111110000100101001001000111101000100101001;
		12'b001101001111: color_data = 108'b000100101001000100101001001000111101000100101001000100101001000100111010001000111101000100101001001000111101;
		12'b001101010000: color_data = 108'b001000111101000100101001001101011111001000111101001000111101000100101001001001001111000100101001001101011111;
		12'b001101010001: color_data = 108'b001101011111001000111101010001111111001001001111001101011111001000111101001101011111001000111101011010001111;
		12'b001101010010: color_data = 108'b010001111111001101011111100010101111001101011111011010001111001001001111010001101111001101011111110111011111;
		12'b001101010011: color_data = 108'b100010101111010001111111011110011111010001101111110111011111001101011111010101111111011010001111101010111111;
		12'b001101010100: color_data = 108'b011110011111100010101111010101111111010101111111101010111111010001101111010001111111110111011111010101111111;
		12'b001101010101: color_data = 108'b010101111111011110011111001101101111010001111111010101111111010101111111001101101111101010111111001101101111;
		12'b001101010110: color_data = 108'b001101101111010101111111001101101111001101101111001101101111010001111111010001101111010101111111001101101111;
		12'b001101010111: color_data = 108'b001101101111001101101111010001111111010001101111001101101111001101101111001101101111001101101111011110001110;
		12'b001101011000: color_data = 108'b010001111111001101101111011110001110001101101111011110001110010001101111010001101111001101101111110011001101;
		12'b001101011001: color_data = 108'b011110001110010001111111110011001110010001101111110011001101001101101111100010011110011110001110111111111111;
		12'b001101011010: color_data = 108'b110011001110011110001110110111011110100010011110111111111111010001101111100110011101110011001101111111111111;
		12'b001101011011: color_data = 108'b110111011110110011001110101110111110100110011101111111111111100010011110011110001110111111111111111011101110;
		12'b001101011100: color_data = 108'b101110111110110111011110011110001111011110001110111011101110100110011101010101111111111111111111101110111101;
		12'b001101011101: color_data = 108'b011110001111101110111110010001111111010101111111101110111101011110001110010001101111111011101110011001111110;
		12'b001101011110: color_data = 108'b010001111111011110001111010001111111010001101111011001111110010101111111010101111111101110111101010001101111;
		12'b001101011111: color_data = 108'b010001111111010001111111010001101111010101111111010001101111010001101111010001111111011001111110001101101111;
		12'b001101100000: color_data = 108'b010001101111010001111111001101101111010001111111001101101111010101111111001101101111010001101111001101101111;
		12'b001101100001: color_data = 108'b001101101111010001101111001101101111001101101111001101101111010001111111001101011111001101101111001101101111;
		12'b001101100010: color_data = 108'b001101101111001101101111001101011111001101011111001101101111001101101111010001101111001101101111010001101111;
		12'b001101100011: color_data = 108'b001101011111001101101111011001111111010001101111010001101111001101011111100010011111001101101111100010011110;
		12'b001101100100: color_data = 108'b011001111111001101011111111011101111100010011111100010011110010001101111111011101111010001101111111011101111;
		12'b001101100101: color_data = 108'b111011101111011001111111111111111111111011101111111011101111100010011111111111111111100010011110111111111111;
		12'b001101100110: color_data = 108'b111111111111111011101111111111111111111111111111111111111111111011101111111111111111111011101111111111111111;
		12'b001101100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110000100: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111100110101111;
		12'b001110000101: color_data = 108'b111011101111111111111111101110111111111111111111100110101111111111111111111011101111111111111111001101011111;
		12'b001110000110: color_data = 108'b101110111111111011101111001101001111111011101111001101011111111111111111101010111111100110101111001001001111;
		12'b001110000111: color_data = 108'b001101001111101110111111001001001111101010111111001001001111111011101111010001011111001101011111000100111011;
		12'b001110001000: color_data = 108'b001001001111001101001111001001001111010001011111000100111011101010111111001001001111001001001111000100101001;
		12'b001110001001: color_data = 108'b001001001111001001001111001001001111001001001111000100101001010001011111001001001111000100111011000100101001;
		12'b001110001010: color_data = 108'b001001001111001001001111001001001111001001001111000100101001001001001111001001001111000100101001000100101010;
		12'b001110001011: color_data = 108'b001001001111001001001111001001001111001001001111000100101010001001001111001001001111000100101001001000111110;
		12'b001110001100: color_data = 108'b001001001111001001001111001000111101001001001111001000111110001001001111001000111101000100101010001000111101;
		12'b001110001101: color_data = 108'b001000111101001001001111000100101001001000111101001000111101001001001111000100101001001000111110000100101001;
		12'b001110001110: color_data = 108'b000100101001001000111101000100101001000100101001000100101001001000111101000100101001001000111101000100101001;
		12'b001110001111: color_data = 108'b000100101001000100101001001000111101000100101001000100101001000100101001001000111101000100101001001000111101;
		12'b001110010000: color_data = 108'b001000111101000100101001001101011111001000111101001000111101000100101001001101011111000100101001001101011111;
		12'b001110010001: color_data = 108'b001101011111001000111101011010001111001101011111001101011111001000111101010001111111001000111101010001101111;
		12'b001110010010: color_data = 108'b011010001111001101011111110111011111010001111111010001101111001101011111100010101111001101011111011010001111;
		12'b001110010011: color_data = 108'b110111011111011010001111101010111111100010101111011010001111010001111111011110011111010001101111011010001111;
		12'b001110010100: color_data = 108'b101010111111110111011111010101111111011110011111011010001111100010101111010101111111011010001111010101111111;
		12'b001110010101: color_data = 108'b010101111111101010111111001101101111010101111111010101111111011110011111001101101111011010001111001101101111;
		12'b001110010110: color_data = 108'b001101101111010101111111001101101111001101101111001101101111010101111111001101101111010101111111001101101111;
		12'b001110010111: color_data = 108'b001101101111001101101111011110001110001101101111001101101111001101101111010001111111001101101111100010101111;
		12'b001110011000: color_data = 108'b011110001110001101101111110011001101010001111111100010101111001101101111011110001110001101101111111111111111;
		12'b001110011001: color_data = 108'b110011001101011110001110111111111111011110001110111111111111010001111111110011001110100010101111111111111111;
		12'b001110011010: color_data = 108'b111111111111110011001101111111111111110011001110111111111111011110001110110111011110111111111111111111111111;
		12'b001110011011: color_data = 108'b111111111111111111111111111011101110110111011110111111111111110011001110101110111110111111111111111111111111;
		12'b001110011100: color_data = 108'b111011101110111111111111101110111101101110111110111111111111110111011110011110001111111111111111110111011110;
		12'b001110011101: color_data = 108'b101110111101111011101110011001111110011110001111110111011110101110111110010001111111111111111111010001000101;
		12'b001110011110: color_data = 108'b011001111110101110111101010001101111010001111111010001000101011110001111010001111111110111011110001000111011;
		12'b001110011111: color_data = 108'b010001101111011001111110001101101111010001111111001000111011010001111111010001101111010001000101001101011111;
		12'b001110100000: color_data = 108'b001101101111010001101111001101101111010001101111001101011111010001111111001101101111001000111011001101101111;
		12'b001110100001: color_data = 108'b001101101111001101101111001101101111001101101111001101101111010001101111001101101111001101011111001101101111;
		12'b001110100010: color_data = 108'b001101101111001101101111010001101111001101101111001101101111001101101111001101011111001101101111001001001001;
		12'b001110100011: color_data = 108'b010001101111001101101111100010011110001101011111001001001001001101101111011001111111001101101111010101010110;
		12'b001110100100: color_data = 108'b100010011110010001101111111011101111011001111111010101010110001101011111111011101111001001001001111011101110;
		12'b001110100101: color_data = 108'b111011101111100010011110111111111111111011101111111011101110011001111111111111111111010101010110111111111111;
		12'b001110100110: color_data = 108'b111111111111111011101111111111111111111111111111111111111111111011101111111111111111111011101110111111111111;
		12'b001110100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b001111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110;
		12'b001111000011: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111100010001100;
		12'b001111000100: color_data = 108'b111111111111111111111111100110101111111111111111100010001100111111111111111011101111111011101110001101001011;
		12'b001111000101: color_data = 108'b100110101111111111111111001101011111111011101111001101001011111111111111101110111111100010001100000100101011;
		12'b001111000110: color_data = 108'b001101011111100110101111001001001111101110111111000100101011111011101111001101001111001101001011000100101011;
		12'b001111000111: color_data = 108'b001001001111001101011111000100111011001101001111000100101011101110111111001001001111000100101011000100101001;
		12'b001111001000: color_data = 108'b000100111011001001001111000100101001001001001111000100101001001101001111001001001111000100101011000100101000;
		12'b001111001001: color_data = 108'b000100101001000100111011000100101001001001001111000100101000001001001111001001001111000100101001000100101000;
		12'b001111001010: color_data = 108'b000100101001000100101001000100101010001001001111000100101000001001001111001001001111000100101000000100101001;
		12'b001111001011: color_data = 108'b000100101010000100101001001000111110001001001111000100101001001001001111001001001111000100101000000100111010;
		12'b001111001100: color_data = 108'b001000111110000100101010001000111101001001001111000100111010001001001111001000111101000100101001000100101010;
		12'b001111001101: color_data = 108'b001000111101001000111110000100101001001000111101000100101010001001001111000100101001000100111010000100101001;
		12'b001111001110: color_data = 108'b000100101001001000111101000100101001000100101001000100101001001000111101000100101001000100101010000100101001;
		12'b001111001111: color_data = 108'b000100101001000100101001001000111101000100101001000100101001000100101001001000111101000100101001000100101010;
		12'b001111010000: color_data = 108'b001000111101000100101001001101011111001000111101000100101010000100101001001101011111000100101001001000111101;
		12'b001111010001: color_data = 108'b001101011111001000111101010001101111001101011111001000111101001000111101011010001111000100101010001101011111;
		12'b001111010010: color_data = 108'b010001101111001101011111011010001111011010001111001101011111001101011111110111011111001000111101010001101111;
		12'b001111010011: color_data = 108'b011010001111010001101111011010001111110111011111010001101111011010001111101010111111001101011111010001101111;
		12'b001111010100: color_data = 108'b011010001111011010001111010101111111101010111111010001101111110111011111010101111111010001101111010001101111;
		12'b001111010101: color_data = 108'b010101111111011010001111001101101111010101111111010001101111101010111111001101101111010001101111001101101111;
		12'b001111010110: color_data = 108'b001101101111010101111111001101101111001101101111001101101111010101111111001101101111010001101111001101101111;
		12'b001111010111: color_data = 108'b001101101111001101101111100010101111001101101111001101101111001101101111011110001110001101101111100110101111;
		12'b001111011000: color_data = 108'b100010101111001101101111111111111111011110001110100110101111001101101111110011001101001101101111111111111111;
		12'b001111011001: color_data = 108'b111111111111100010101111111111111111110011001101111111111111011110001110111111111111100110101111111111111111;
		12'b001111011010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111110011001101111111111111111111111111111111111111;
		12'b001111011011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111;
		12'b001111011100: color_data = 108'b111111111111111111111111110111011110111011101110111111111111111111111111101110111101111111111111111011101110;
		12'b001111011101: color_data = 108'b110111011110111111111111010001000101101110111101111011101110111011101110011001111110111111111111001100110011;
		12'b001111011110: color_data = 108'b010001000101110111011110001000111011011001111110001100110011101110111101010001101111111011101110001000100101;
		12'b001111011111: color_data = 108'b001000111011010001000101001101011111010001101111001000100101011001111110001101101111001100110011001000111010;
		12'b001111100000: color_data = 108'b001101011111001000111011001101101111001101101111001000111010010001101111001101101111001000100101001001011111;
		12'b001111100001: color_data = 108'b001101101111001101011111001101101111001101101111001001011111001101101111001101101111001000111010001101101111;
		12'b001111100010: color_data = 108'b001101101111001101101111001001001001001101101111001101101111001101101111010001101111001001011111001000111000;
		12'b001111100011: color_data = 108'b001001001001001101101111010101010110010001101111001000111000001101101111100010011110001101101111010101010101;
		12'b001111100100: color_data = 108'b010101010110001001001001111011101110100010011110010101010101010001101111111011101111001000111000111011101110;
		12'b001111100101: color_data = 108'b111011101110010101010110111111111111111011101111111011101110100010011110111111111111010101010101111111111111;
		12'b001111100110: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111011101111111111111111111011101110111111111111;
		12'b001111100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b001111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000000010: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111111111111111111111111111011101110;
		12'b010000000011: color_data = 108'b111011101110111111111111100010001100111111111111111011101110111111111111111111111111111111111111011101111011;
		12'b010000000100: color_data = 108'b100010001100111011101110001101001011111111111111011101111011111111111111100110101111111011101110010101101010;
		12'b010000000101: color_data = 108'b001101001011100010001100000100101011100110101111010101101010111111111111001101011111011101111011010101101010;
		12'b010000000110: color_data = 108'b000100101011001101001011000100101011001101011111010101101010100110101111001001001111010101101010010101101010;
		12'b010000000111: color_data = 108'b000100101011000100101011000100101001001001001111010101101010001101011111000100111011010101101010010101101010;
		12'b010000001000: color_data = 108'b000100101001000100101011000100101000000100111011010101101010001001001111000100101001010101101010010101101010;
		12'b010000001001: color_data = 108'b000100101000000100101001000100101000000100101001010101101010000100111011000100101001010101101010010001011010;
		12'b010000001010: color_data = 108'b000100101000000100101000000100101001000100101001010001011010000100101001000100101010010101101010000100101001;
		12'b010000001011: color_data = 108'b000100101001000100101000000100111010000100101010000100101001000100101001001000111110010001011010000100101000;
		12'b010000001100: color_data = 108'b000100111010000100101001000100101010001000111110000100101000000100101010001000111101000100101001000100101000;
		12'b010000001101: color_data = 108'b000100101010000100111010000100101001001000111101000100101000001000111110000100101001000100101000000100101001;
		12'b010000001110: color_data = 108'b000100101001000100101010000100101001000100101001000100101001001000111101000100101001000100101000000100101001;
		12'b010000001111: color_data = 108'b000100101001000100101001000100101010000100101001000100101001000100101001001000111101000100101001000100101000;
		12'b010000010000: color_data = 108'b000100101010000100101001001000111101001000111101000100101000000100101001001101011111000100101001000100111011;
		12'b010000010001: color_data = 108'b001000111101000100101010001101011111001101011111000100111011001000111101010001101111000100101000001001001111;
		12'b010000010010: color_data = 108'b001101011111001000111101010001101111010001101111001001001111001101011111011010001111000100111011001101011111;
		12'b010000010011: color_data = 108'b010001101111001101011111010001101111011010001111001101011111010001101111011010001111001001001111001101011111;
		12'b010000010100: color_data = 108'b010001101111010001101111010001101111011010001111001101011111011010001111010101111111001101011111001101011111;
		12'b010000010101: color_data = 108'b010001101111010001101111001101101111010101111111001101011111011010001111001101101111001101011111001101011111;
		12'b010000010110: color_data = 108'b001101101111010001101111001101101111001101101111001101011111010101111111001101101111001101011111001101011111;
		12'b010000010111: color_data = 108'b001101101111001101101111100110101111001101101111001101011111001101101111100010101111001101011111100110101111;
		12'b010000011000: color_data = 108'b100110101111001101101111111111111111100010101111100110101111001101101111111111111111001101011111111111111111;
		12'b010000011001: color_data = 108'b111111111111100110101111111111111111111111111111111111111111100010101111111111111111100110101111111111111111;
		12'b010000011010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000011011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000011100: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111110111011110111111111111111011101110;
		12'b010000011101: color_data = 108'b111011101110111111111111001100110011110111011110111011101110111111111111010001000101111111111111001100110011;
		12'b010000011110: color_data = 108'b001100110011111011101110001000100101010001000101001100110011110111011110001000111011111011101110001000100001;
		12'b010000011111: color_data = 108'b001000100101001100110011001000111010001000111011001000100001010001000101001101011111001100110011001000110110;
		12'b010000100000: color_data = 108'b001000111010001000100101001001011111001101011111001000110110001000111011001101101111001000100001001101011111;
		12'b010000100001: color_data = 108'b001001011111001000111010001101101111001101101111001101011111001101011111001101101111001000110110001101011100;
		12'b010000100010: color_data = 108'b001101101111001001011111001000111000001101101111001101011100001101101111001001001001001101011111001000110110;
		12'b010000100011: color_data = 108'b001000111000001101101111010101010101001001001001001000110110001101101111010101010110001101011100010101010101;
		12'b010000100100: color_data = 108'b010101010101001000111000111011101110010101010110010101010101001001001001111011101110001000110110111011101110;
		12'b010000100101: color_data = 108'b111011101110010101010101111111111111111011101110111011101110010101010110111111111111010101010101111111111111;
		12'b010000100110: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111011101110111111111111111011101110111111111111;
		12'b010000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001000010: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111011101110111111111111111111111111;
		12'b010001000011: color_data = 108'b111011101110111111111111011101111011111011101110111111111111111111111111100010001100111111111111111011101111;
		12'b010001000100: color_data = 108'b011101111011111011101110010101101010100010001100111011101111111011101110001101001011111111111111111011101111;
		12'b010001000101: color_data = 108'b010101101010011101111011010101101010001101001011111011101111100010001100000100101011111011101111111011101111;
		12'b010001000110: color_data = 108'b010101101010010101101010010101101010000100101011111011101111001101001011000100101011111011101111111011101111;
		12'b010001000111: color_data = 108'b010101101010010101101010010101101010000100101011111011101111000100101011000100101001111011101111111011101111;
		12'b010001001000: color_data = 108'b010101101010010101101010010101101010000100101001111011101111000100101011000100101000111011101111111111111111;
		12'b010001001001: color_data = 108'b010101101010010101101010010001011010000100101000111111111111000100101001000100101000111011101111110011001110;
		12'b010001001010: color_data = 108'b010001011010010101101010000100101001000100101000110011001110000100101000000100101001111111111111001101001001;
		12'b010001001011: color_data = 108'b000100101001010001011010000100101000000100101001001101001001000100101000000100111010110011001110001000111001;
		12'b010001001100: color_data = 108'b000100101000000100101001000100101000000100111010001000111001000100101001000100101010001101001001001000111001;
		12'b010001001101: color_data = 108'b000100101000000100101000000100101001000100101010001000111001000100111010000100101001001000111001000100101001;
		12'b010001001110: color_data = 108'b000100101001000100101000000100101001000100101001000100101001000100101010000100101001001000111001000100101001;
		12'b010001001111: color_data = 108'b000100101001000100101001000100101000000100101001000100101001000100101001000100101010000100101001000100101000;
		12'b010001010000: color_data = 108'b000100101000000100101001000100111011000100101010000100101000000100101001001000111101000100101001000100111011;
		12'b010001010001: color_data = 108'b000100111011000100101000001001001111001000111101000100111011000100101010001101011111000100101000001001001111;
		12'b010001010010: color_data = 108'b001001001111000100111011001101011111001101011111001001001111001000111101010001101111000100111011001001001111;
		12'b010001010011: color_data = 108'b001101011111001001001111001101011111010001101111001001001111001101011111010001101111001001001111001001001111;
		12'b010001010100: color_data = 108'b001101011111001101011111001101011111010001101111001001001111010001101111010001101111001001001111001001001111;
		12'b010001010101: color_data = 108'b001101011111001101011111001101011111010001101111001001001111010001101111001101101111001001001111001001001111;
		12'b010001010110: color_data = 108'b001101011111001101011111001101011111001101101111001001001111010001101111001101101111001001001111001101011111;
		12'b010001010111: color_data = 108'b001101011111001101011111100110101111001101101111001101011111001101101111100110101111001001001111100010101111;
		12'b010001011000: color_data = 108'b100110101111001101011111111111111111100110101111100010101111001101101111111111111111001101011111111111111111;
		12'b010001011001: color_data = 108'b111111111111100110101111111111111111111111111111111111111111100110101111111111111111100010101111111111111111;
		12'b010001011010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001011011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001011100: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111011101110111111111111111011101110;
		12'b010001011101: color_data = 108'b111011101110111111111111001100110011111011101110111011101110111111111111001100110011111111111111001100110011;
		12'b010001011110: color_data = 108'b001100110011111011101110001000100001001100110011001100110011111011101110001000100101111011101110001000100010;
		12'b010001011111: color_data = 108'b001000100001001100110011001000110110001000100101001000100010001100110011001000111010001100110011001101000110;
		12'b010001100000: color_data = 108'b001000110110001000100001001101011111001000111010001101000110001000100101001001011111001000100010011001111110;
		12'b010001100001: color_data = 108'b001101011111001000110110001101011100001001011111011001111110001000111010001101101111001101000110001100110101;
		12'b010001100010: color_data = 108'b001101011100001101011111001000110110001101101111001100110101001001011111001000111000011001111110001000100010;
		12'b010001100011: color_data = 108'b001000110110001101011100010101010101001000111000001000100010001101101111010101010101001100110101010101010101;
		12'b010001100100: color_data = 108'b010101010101001000110110111011101110010101010101010101010101001000111000111011101110001000100010111011101110;
		12'b010001100101: color_data = 108'b111011101110010101010101111111111111111011101110111011101110010101010101111111111111010101010101111111111111;
		12'b010001100110: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111011101110111111111111111011101110111111111111;
		12'b010001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111;
		12'b010010000011: color_data = 108'b111111111111111111111111111011101111111011101110111111111111111111111111011101111011111111111111111111111111;
		12'b010010000100: color_data = 108'b111011101111111111111111111011101111011101111011111111111111111011101110010101101010111111111111111111111111;
		12'b010010000101: color_data = 108'b111011101111111011101111111011101111010101101010111111111111011101111011010101101010111111111111111111111111;
		12'b010010000110: color_data = 108'b111011101111111011101111111011101111010101101010111111111111010101101010010101101010111111111111111111111111;
		12'b010010000111: color_data = 108'b111011101111111011101111111011101111010101101010111111111111010101101010010101101010111111111111111111111111;
		12'b010010001000: color_data = 108'b111011101111111011101111111111111111010101101010111111111111010101101010010101101010111111111111111111111111;
		12'b010010001001: color_data = 108'b111111111111111011101111110011001110010101101010111111111111010101101010010001011010111111111111111011101111;
		12'b010010001010: color_data = 108'b110011001110111111111111001101001001010001011010111011101111010101101010000100101001111111111111110011001110;
		12'b010010001011: color_data = 108'b001101001001110011001110001000111001000100101001110011001110010001011010000100101000111011101111110011011110;
		12'b010010001100: color_data = 108'b001000111001001101001001001000111001000100101000110011011110000100101001000100101000110011001110100010001100;
		12'b010010001101: color_data = 108'b001000111001001000111001000100101001000100101000100010001100000100101000000100101001110011011110000100101001;
		12'b010010001110: color_data = 108'b000100101001001000111001000100101001000100101001000100101001000100101000000100101001100010001100000100101001;
		12'b010010001111: color_data = 108'b000100101001000100101001000100101000000100101001000100101001000100101001000100101000000100101001000100101001;
		12'b010010010000: color_data = 108'b000100101000000100101001000100111011000100101000000100101001000100101001000100111011000100101001000100101001;
		12'b010010010001: color_data = 108'b000100111011000100101000001001001111000100111011000100101001000100101000001001001111000100101001000100101010;
		12'b010010010010: color_data = 108'b001001001111000100111011001001001111001001001111000100101010000100111011001101011111000100101001001001001111;
		12'b010010010011: color_data = 108'b001001001111001001001111001001001111001101011111001001001111001001001111001101011111000100101010001001001111;
		12'b010010010100: color_data = 108'b001001001111001001001111001001001111001101011111001001001111001101011111001101011111001001001111001001001111;
		12'b010010010101: color_data = 108'b001001001111001001001111001001001111001101011111001001001111001101011111001101011111001001001111001001001111;
		12'b010010010110: color_data = 108'b001001001111001001001111001101011111001101011111001001001111001101011111001101011111001001001111001001001111;
		12'b010010010111: color_data = 108'b001101011111001001001111100010101111001101011111001001001111001101011111100110101111001001001111010001101111;
		12'b010010011000: color_data = 108'b100010101111001101011111111111111111100110101111010001101111001101011111111111111111001001001111100110101111;
		12'b010010011001: color_data = 108'b111111111111100010101111111111111111111111111111100110101111100110101111111111111111010001101111111111111111;
		12'b010010011010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110101111111111111111;
		12'b010010011011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010011100: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111011101110111111111111111011101110;
		12'b010010011101: color_data = 108'b111011101110111111111111001100110011111011101110111011101110111111111111001100110011111111111111001100110011;
		12'b010010011110: color_data = 108'b001100110011111011101110001000100010001100110011001100110011111011101110001000100001111011101110000100010001;
		12'b010010011111: color_data = 108'b001000100010001100110011001101000110001000100001000100010001001100110011001000110110001100110011010101010110;
		12'b010010100000: color_data = 108'b001101000110001000100010011001111110001000110110010101010110001000100001001101011111000100010001110111011110;
		12'b010010100001: color_data = 108'b011001111110001101000110001100110101001101011111110111011110001000110110001101011100010101010110010001000100;
		12'b010010100010: color_data = 108'b001100110101011001111110001000100010001101011100010001000100001101011111001000110110110111011110010001000101;
		12'b010010100011: color_data = 108'b001000100010001100110101010101010101001000110110010001000101001101011100010101010101010001000100100010001001;
		12'b010010100100: color_data = 108'b010101010101001000100010111011101110010101010101100010001001001000110110111011101110010001000101111011101110;
		12'b010010100101: color_data = 108'b111011101110010101010101111111111111111011101110111011101110010101010101111111111111100010001001111111111111;
		12'b010010100110: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111011101110111111111111111011101110111111111111;
		12'b010010100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111;
		12'b010011000100: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111111111111111011101111111111111111111111111111;
		12'b010011000101: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111011101111111011101111111111111111111111111111;
		12'b010011000110: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111011101111111011101111111111111111111111111111;
		12'b010011000111: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111011101111111011101111111111111111111111111111;
		12'b010011001000: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111011101111111111111111111111111111111111111111;
		12'b010011001001: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111011101111110011001110111111111111111111111111;
		12'b010011001010: color_data = 108'b111011101111111111111111110011001110110011001110111111111111111111111111001101001001111111111111111111111111;
		12'b010011001011: color_data = 108'b110011001110111011101111110011011110001101001001111111111111110011001110001000111001111111111111101010111111;
		12'b010011001100: color_data = 108'b110011011110110011001110100010001100001000111001101010111111001101001001001000111001111111111111011001111110;
		12'b010011001101: color_data = 108'b100010001100110011011110000100101001001000111001011001111110001000111001000100101001101010111111001000111100;
		12'b010011001110: color_data = 108'b000100101001100010001100000100101001000100101001001000111100001000111001000100101001011001111110000100101001;
		12'b010011001111: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101000001000111100000100101001;
		12'b010011010000: color_data = 108'b000100101001000100101001000100101001000100101000000100101001000100101001000100111011000100101001000100101001;
		12'b010011010001: color_data = 108'b000100101001000100101001000100101010000100111011000100101001000100101000001001001111000100101001000100101001;
		12'b010011010010: color_data = 108'b000100101010000100101001001001001111001001001111000100101001000100111011001001001111000100101001000100111011;
		12'b010011010011: color_data = 108'b001001001111000100101010001001001111001001001111000100111011001001001111001001001111000100101001001000111110;
		12'b010011010100: color_data = 108'b001001001111001001001111001001001111001001001111001000111110001001001111001001001111000100111011001101001110;
		12'b010011010101: color_data = 108'b001001001111001001001111001001001111001001001111001101001110001001001111001001001111001000111110011101101010;
		12'b010011010110: color_data = 108'b001001001111001001001111001001001111001001001111011101101010001001001111001101011111001101001110100110011110;
		12'b010011010111: color_data = 108'b001001001111001001001111010001101111001101011111100110011110001001001111100010101111011101101010101010111111;
		12'b010011011000: color_data = 108'b010001101111001001001111100110101111100010101111101010111111001101011111111111111111100110011110101110111111;
		12'b010011011001: color_data = 108'b100110101111010001101111111111111111111111111111101110111111100010101111111111111111101010111111101010111111;
		12'b010011011010: color_data = 108'b111111111111100110101111111111111111111111111111101010111111111111111111111111111111101110111111111011101111;
		12'b010011011011: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111101010111111111111111111;
		12'b010011011100: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111011101110111011101111111111111111;
		12'b010011011101: color_data = 108'b111011101110111111111111001100110011111011101110111111111111111111111111001100110011111111111111101010101010;
		12'b010011011110: color_data = 108'b001100110011111011101110000100010001001100110011101010101010111011101110001000100010111111111111100110011001;
		12'b010011011111: color_data = 108'b000100010001001100110011010101010110001000100010100110011001001100110011001101000110101010101010101010101001;
		12'b010011100000: color_data = 108'b010101010110000100010001110111011110001101000110101010101001001000100010011001111110100110011001110010111001;
		12'b010011100001: color_data = 108'b110111011110010101010110010001000100011001111110110010111001001101000110001100110101101010101001011001100110;
		12'b010011100010: color_data = 108'b010001000100110111011110010001000101001100110101011001100110011001111110001000100010110010111001010101010101;
		12'b010011100011: color_data = 108'b010001000101010001000100100010001001001000100010010101010101001100110101010101010101011001100110011001100111;
		12'b010011100100: color_data = 108'b100010001001010001000101111011101110010101010101011001100111001000100010111011101110010101010101101110111011;
		12'b010011100101: color_data = 108'b111011101110100010001001111111111111111011101110101110111011010101010101111111111111011001100111111011101110;
		12'b010011100110: color_data = 108'b111111111111111011101110111111111111111111111111111011101110111011101110111111111111101110111011111111111111;
		12'b010011100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111;
		12'b010011101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111;
		12'b010100001001: color_data = 108'b111111111111111111111111111111111111111111111111110111101111111111111111111011101111111111111111110011001111;
		12'b010100001010: color_data = 108'b111111111111111111111111111111111111111011101111110011001111111111111111110011001110110111101111110011001111;
		12'b010100001011: color_data = 108'b111111111111111111111111101010111111110011001110110011001111111011101111110011011110110011001111010101101111;
		12'b010100001100: color_data = 108'b101010111111111111111111011001111110110011011110010101101111110011001110100010001100110011001111001001001111;
		12'b010100001101: color_data = 108'b011001111110101010111111001000111100100010001100001001001111110011011110000100101001010101101111001001001111;
		12'b010100001110: color_data = 108'b001000111100011001111110000100101001000100101001001001001111100010001100000100101001001001001111000100101001;
		12'b010100001111: color_data = 108'b000100101001001000111100000100101001000100101001000100101001000100101001000100101001001001001111000100101001;
		12'b010100010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010100010001: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101010000100101001000100101001;
		12'b010100010010: color_data = 108'b000100101001000100101001000100111011000100101010000100101001000100101001001001001111000100101001000100101000;
		12'b010100010011: color_data = 108'b000100111011000100101001001000111110001001001111000100101000000100101010001001001111000100101001001100111011;
		12'b010100010100: color_data = 108'b001000111110000100111011001101001110001001001111001100111011001001001111001001001111000100101000011001101011;
		12'b010100010101: color_data = 108'b001101001110001000111110011101101010001001001111011001101011001001001111001001001111001100111011110010010110;
		12'b010100010110: color_data = 108'b011101101010001101001110100110011110001001001111110010010110001001001111001001001111011001101011111111011100;
		12'b010100010111: color_data = 108'b100110011110011101101010101010111111001001001111111111011100001001001111010001101111110010010110111111111110;
		12'b010100011000: color_data = 108'b101010111111100110011110101110111111010001101111111111111110001001001111100110101111111111011100111011101110;
		12'b010100011001: color_data = 108'b101110111111101010111111101010111111100110101111111011101110010001101111111111111111111111111110100010101111;
		12'b010100011010: color_data = 108'b101010111111101110111111111011101111111111111111100010101111100110101111111111111111111011101110110111011111;
		12'b010100011011: color_data = 108'b111011101111101010111111111111111111111111111111110111011111111111111111111111111111100010101111111111111111;
		12'b010100011100: color_data = 108'b111111111111111011101111111111111111111111111111111111111111111111111111111011101110110111011111111111111111;
		12'b010100011101: color_data = 108'b111111111111111111111111101010101010111011101110111111111111111111111111001100110011111111111111111111111111;
		12'b010100011110: color_data = 108'b101010101010111111111111100110011001001100110011111111111111111011101110000100010001111111111111111111111111;
		12'b010100011111: color_data = 108'b100110011001101010101010101010101001000100010001111111111111001100110011010101010110111111111111111111011100;
		12'b010100100000: color_data = 108'b101010101001100110011001110010111001010101010110111111011100000100010001110111011110111111111111110010000110;
		12'b010100100001: color_data = 108'b110010111001101010101001011001100110110111011110110010000110010101010110010001000100111111011100011101110111;
		12'b010100100010: color_data = 108'b011001100110110010111001010101010101010001000100011101110111110111011110010001000101110010000110010001000100;
		12'b010100100011: color_data = 108'b010101010101011001100110011001100111010001000101010001000100010001000100100010001001011101110111001100110011;
		12'b010100100100: color_data = 108'b011001100111010101010101101110111011100010001001001100110011010001000101111011101110010001000100011001100111;
		12'b010100100101: color_data = 108'b101110111011011001100111111011101110111011101110011001100111100010001001111111111111001100110011110111011101;
		12'b010100100110: color_data = 108'b111011101110101110111011111111111111111111111111110111011101111011101110111111111111011001100111111111111111;
		12'b010100100111: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111111111111111111111111110111011101111111111111;
		12'b010100101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101001000: color_data = 108'b111111111111111111111111110111101111111111111111111111111111111111111111111111111111111111111111100110101111;
		12'b010101001001: color_data = 108'b110111101111111111111111110011001111111111111111100110101111111111111111111111111111111111111111001101001111;
		12'b010101001010: color_data = 108'b110011001111110111101111110011001111111111111111001101001111111111111111111111111111100110101111001101001111;
		12'b010101001011: color_data = 108'b110011001111110011001111010101101111111111111111001101001111111111111111101010111111001101001111001001001111;
		12'b010101001100: color_data = 108'b010101101111110011001111001001001111101010111111001001001111111111111111011001111110001101001111001001001111;
		12'b010101001101: color_data = 108'b001001001111010101101111001001001111011001111110001001001111101010111111001000111100001001001111001001001110;
		12'b010101001110: color_data = 108'b001001001111001001001111000100101001001000111100001001001110011001111110000100101001001001001111000100101001;
		12'b010101001111: color_data = 108'b000100101001001001001111000100101001000100101001000100101001001000111100000100101001001001001110000100101001;
		12'b010101010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010101010001: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010101010010: color_data = 108'b000100101001000100101001000100101000000100101001000100101001000100101001000100111011000100101001000100101001;
		12'b010101010011: color_data = 108'b000100101000000100101001001100111011000100111011000100101001000100101001001000111110000100101001011001010111;
		12'b010101010100: color_data = 108'b001100111011000100101000011001101011001000111110011001010111000100111011001101001110000100101001110010000110;
		12'b010101010101: color_data = 108'b011001101011001100111011110010010110001101001110110010000110001000111110011101101010011001010111111110111001;
		12'b010101010110: color_data = 108'b110010010110011001101011111111011100011101101010111110111001001101001110100110011110110010000110111111001010;
		12'b010101010111: color_data = 108'b111111011100110010010110111111111110100110011110111111001010011101101010101010111111111110111001111111001010;
		12'b010101011000: color_data = 108'b111111111110111111011100111011101110101010111111111111001010100110011110101110111111111111001010111111001011;
		12'b010101011001: color_data = 108'b111011101110111111111110100010101111101110111111111111001011101010111111101010111111111111001010111111111111;
		12'b010101011010: color_data = 108'b100010101111111011101110110111011111101010111111111111111111101110111111111011101111111111001011111111111111;
		12'b010101011011: color_data = 108'b110111011111100010101111111111111111111011101111111111111111101010111111111111111111111111111111111111111111;
		12'b010101011100: color_data = 108'b111111111111110111011111111111111111111111111111111111111111111011101111111111111111111111111111111111111111;
		12'b010101011101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111101010101010111111111111111111111111;
		12'b010101011110: color_data = 108'b111111111111111111111111111111111111101010101010111111111111111111111111100110011001111111111111111111011100;
		12'b010101011111: color_data = 108'b111111111111111111111111111111011100100110011001111111011100101010101010101010101001111111111111111111001010;
		12'b010101100000: color_data = 108'b111111011100111111111111110010000110101010101001111111001010100110011001110010111001111111011100111010111001;
		12'b010101100001: color_data = 108'b110010000110111111011100011101110111110010111001111010111001101010101001011001100110111111001010010101000100;
		12'b010101100010: color_data = 108'b011101110111110010000110010001000100011001100110010101000100110010111001010101010101111010111001001000100010;
		12'b010101100011: color_data = 108'b010001000100011101110111001100110011010101010101001000100010011001100110011001100111010101000100001000100010;
		12'b010101100100: color_data = 108'b001100110011010001000100011001100111011001100111001000100010010101010101101110111011001000100010001100110011;
		12'b010101100101: color_data = 108'b011001100111001100110011110111011101101110111011001100110011011001100111111011101110001000100010110011001100;
		12'b010101100110: color_data = 108'b110111011101011001100111111111111111111011101110110011001100101110111011111111111111001100110011111111111111;
		12'b010101100111: color_data = 108'b111111111111110111011101111111111111111111111111111111111111111011101110111111111111110011001100111111111111;
		12'b010101101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b010110000111: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111100010011111;
		12'b010110001000: color_data = 108'b111111111111111111111111100110101111111111111111100010011111111111111111110111101111111011101111010001011111;
		12'b010110001001: color_data = 108'b100110101111111111111111001101001111110111101111010001011111111111111111110011001111100010011111001001001111;
		12'b010110001010: color_data = 108'b001101001111100110101111001101001111110011001111001001001111110111101111110011001111010001011111001001001111;
		12'b010110001011: color_data = 108'b001101001111001101001111001001001111110011001111001001001111110011001111010101101111001001001111001000111100;
		12'b010110001100: color_data = 108'b001001001111001101001111001001001111010101101111001000111100110011001111001001001111001001001111000100101010;
		12'b010110001101: color_data = 108'b001001001111001001001111001001001110001001001111000100101010010101101111001001001111001000111100000100101010;
		12'b010110001110: color_data = 108'b001001001110001001001111000100101001001001001111000100101010001001001111000100101001000100101010000100101001;
		12'b010110001111: color_data = 108'b000100101001001001001110000100101001000100101001000100101001001001001111000100101001000100101010000100101001;
		12'b010110010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010110010001: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010110010010: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101000000100101001000100101001;
		12'b010110010011: color_data = 108'b000100101001000100101001011001010111000100101000000100101001000100101001001100111011000100101001011001010110;
		12'b010110010100: color_data = 108'b011001010111000100101001110010000110001100111011011001010110000100101000011001101011000100101001110010010110;
		12'b010110010101: color_data = 108'b110010000110011001010111111110111001011001101011110010010110001100111011110010010110011001010110111111001001;
		12'b010110010110: color_data = 108'b111110111001110010000110111111001010110010010110111111001001011001101011111111011100110010010110111111001010;
		12'b010110010111: color_data = 108'b111111001010111110111001111111001010111111011100111111001010110010010110111111111110111111001001111111001010;
		12'b010110011000: color_data = 108'b111111001010111111001010111111001011111111111110111111001010111111011100111011101110111111001010111111001010;
		12'b010110011001: color_data = 108'b111111001011111111001010111111111111111011101110111111001010111111111110100010101111111111001010111111011011;
		12'b010110011010: color_data = 108'b111111111111111111001011111111111111100010101111111111011011111011101110110111011111111111001010111111011011;
		12'b010110011011: color_data = 108'b111111111111111111111111111111111111110111011111111111011011100010101111111111111111111111011011111111011011;
		12'b010110011100: color_data = 108'b111111111111111111111111111111111111111111111111111111011011110111011111111111111111111111011011111111011011;
		12'b010110011101: color_data = 108'b111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111011011111111011011;
		12'b010110011110: color_data = 108'b111111111111111111111111111111011100111111111111111111011011111111111111111111111111111111011011111111001010;
		12'b010110011111: color_data = 108'b111111011100111111111111111111001010111111111111111111001010111111111111111111011100111111011011111111001010;
		12'b010110100000: color_data = 108'b111111001010111111011100111010111001111111011100111111001010111111111111110010000110111111001010111111001010;
		12'b010110100001: color_data = 108'b111010111001111111001010010101000100110010000110111111001010111111011100011101110111111111001010110011001011;
		12'b010110100010: color_data = 108'b010101000100111010111001001000100010011101110111110011001011110010000110010001000100111111001010101111001100;
		12'b010110100011: color_data = 108'b001000100010010101000100001000100010010001000100101111001100011101110111001100110011110011001011101110111011;
		12'b010110100100: color_data = 108'b001000100010001000100010001100110011001100110011101110111011010001000100011001100111101111001100110011001100;
		12'b010110100101: color_data = 108'b001100110011001000100010110011001100011001100111110011001100001100110011110111011101101110111011111011101110;
		12'b010110100110: color_data = 108'b110011001100001100110011111111111111110111011101111011101110011001100111111111111111110011001100111111111111;
		12'b010110100111: color_data = 108'b111111111111110011001100111111111111111111111111111111111111110111011101111111111111111011101110111111111111;
		12'b010110101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b010111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111000110: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b010111000111: color_data = 108'b111011101111111111111111100010011111111111111111111011101111111111111111111111111111111111111111010101101111;
		12'b010111001000: color_data = 108'b100010011111111011101111010001011111111111111111010101101111111111111111100110101111111011101111001000111110;
		12'b010111001001: color_data = 108'b010001011111100010011111001001001111100110101111001000111110111111111111001101001111010101101111001000111100;
		12'b010111001010: color_data = 108'b001001001111010001011111001001001111001101001111001000111100100110101111001101001111001000111110001000111100;
		12'b010111001011: color_data = 108'b001001001111001001001111001000111100001101001111001000111100001101001111001001001111001000111100000100101010;
		12'b010111001100: color_data = 108'b001000111100001001001111000100101010001001001111000100101010001101001111001001001111001000111100000100101000;
		12'b010111001101: color_data = 108'b000100101010001000111100000100101010001001001111000100101000001001001111001001001110000100101010000100101001;
		12'b010111001110: color_data = 108'b000100101010000100101010000100101001001001001110000100101001001001001111000100101001000100101000000100101001;
		12'b010111001111: color_data = 108'b000100101001000100101010000100101001000100101001000100101001001001001110000100101001000100101001000100101001;
		12'b010111010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010111010001: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010111010010: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b010111010011: color_data = 108'b000100101001000100101001011001010110000100101001000100101001000100101001011001010111000100101001010001000111;
		12'b010111010100: color_data = 108'b011001010110000100101001110010010110011001010111010001000111000100101001110010000110000100101001100001100111;
		12'b010111010101: color_data = 108'b110010010110011001010110111111001001110010000110100001100111011001010111111110111001010001000111110110101000;
		12'b010111010110: color_data = 108'b111111001001110010010110111111001010111110111001110110101000110010000110111111001010100001100111111110111001;
		12'b010111010111: color_data = 108'b111111001010111111001001111111001010111111001010111110111001111110111001111111001010110110101000111111001010;
		12'b010111011000: color_data = 108'b111111001010111111001010111111001010111111001010111111001010111111001010111111001011111110111001111111001010;
		12'b010111011001: color_data = 108'b111111001010111111001010111111011011111111001011111111001010111111001010111111111111111111001010111111001010;
		12'b010111011010: color_data = 108'b111111011011111111001010111111011011111111111111111111001010111111001011111111111111111111001010111111001010;
		12'b010111011011: color_data = 108'b111111011011111111011011111111011011111111111111111111001010111111111111111111111111111111001010111111001010;
		12'b010111011100: color_data = 108'b111111011011111111011011111111011011111111111111111111001010111111111111111111111111111111001010111111001001;
		12'b010111011101: color_data = 108'b111111011011111111011011111111011011111111111111111111001001111111111111111111111111111111001010111010101000;
		12'b010111011110: color_data = 108'b111111011011111111011011111111001010111111111111111010101000111111111111111111011100111111001001111010101000;
		12'b010111011111: color_data = 108'b111111001010111111011011111111001010111111011100111010101000111111111111111111001010111010101000110110010111;
		12'b010111100000: color_data = 108'b111111001010111111001010111111001010111111001010110110010111111111011100111010111001111010101000110101110110;
		12'b010111100001: color_data = 108'b111111001010111111001010110011001011111010111001110101110110111111001010010101000100110110010111111011011101;
		12'b010111100010: color_data = 108'b110011001011111111001010101111001100010101000100111011011101111010111001001000100010110101110110111111111111;
		12'b010111100011: color_data = 108'b101111001100110011001011101110111011001000100010111111111111010101000100001000100010111011011101111111111111;
		12'b010111100100: color_data = 108'b101110111011101111001100110011001100001000100010111111111111001000100010001100110011111111111111111111111111;
		12'b010111100101: color_data = 108'b110011001100101110111011111011101110001100110011111111111111001000100010110011001100111111111111111111111111;
		12'b010111100110: color_data = 108'b111011101110110011001100111111111111110011001100111111111111001100110011111111111111111111111111111111111111;
		12'b010111100111: color_data = 108'b111111111111111011101110111111111111111111111111111111111111110011001100111111111111111111111111111111111111;
		12'b010111101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b010111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b011000000110: color_data = 108'b111111111111111111111111111011101111111111111111111011101111111111111111111011101111111111111111110011011111;
		12'b011000000111: color_data = 108'b111011101111111111111111010101101111111011101111110011011111111111111111100010011111111011101111010101101110;
		12'b011000001000: color_data = 108'b010101101111111011101111001000111110100010011111010101101110111011101111010001011111110011011111000100111100;
		12'b011000001001: color_data = 108'b001000111110010101101111001000111100010001011111000100111100100010011111001001001111010101101110000100101000;
		12'b011000001010: color_data = 108'b001000111100001000111110001000111100001001001111000100101000010001011111001001001111000100111100000100101001;
		12'b011000001011: color_data = 108'b001000111100001000111100000100101010001001001111000100101001001001001111001000111100000100101000000100101001;
		12'b011000001100: color_data = 108'b000100101010001000111100000100101000001000111100000100101001001001001111000100101010000100101001000100101001;
		12'b011000001101: color_data = 108'b000100101000000100101010000100101001000100101010000100101001001000111100000100101010000100101001000100101001;
		12'b011000001110: color_data = 108'b000100101001000100101000000100101001000100101010000100101001000100101010000100101001000100101001000100101001;
		12'b011000001111: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101010000100101001000100101001000100101001;
		12'b011000010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b011000010001: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b011000010010: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101000;
		12'b011000010011: color_data = 108'b000100101001000100101001010001000111000100101001000100101000000100101001011001010110000100101001000100101000;
		12'b011000010100: color_data = 108'b010001000111000100101001100001100111011001010110000100101000000100101001110010010110000100101000001100111000;
		12'b011000010101: color_data = 108'b100001100111010001000111110110101000110010010110001100111000011001010110111111001001000100101000100101110110;
		12'b011000010110: color_data = 108'b110110101000100001100111111110111001111111001001100101110110110010010110111111001010001100111000110110101000;
		12'b011000010111: color_data = 108'b111110111001110110101000111111001010111111001010110110101000111111001001111111001010100101110110111110111001;
		12'b011000011000: color_data = 108'b111111001010111110111001111111001010111111001010111110111001111111001010111111001010110110101000111110111001;
		12'b011000011001: color_data = 108'b111111001010111111001010111111001010111111001010111110111001111111001010111111011011111110111001111110111001;
		12'b011000011010: color_data = 108'b111111001010111111001010111111001010111111011011111110111001111111001010111111011011111110111001111110111001;
		12'b011000011011: color_data = 108'b111111001010111111001010111111001010111111011011111110111001111111011011111111011011111110111001111110111001;
		12'b011000011100: color_data = 108'b111111001010111111001010111111001001111111011011111110111001111111011011111111011011111110111001111010101000;
		12'b011000011101: color_data = 108'b111111001001111111001010111010101000111111011011111010101000111111011011111111011011111110111001101101110100;
		12'b011000011110: color_data = 108'b111010101000111111001001111010101000111111011011101101110100111111011011111111001010111010101000101001100100;
		12'b011000011111: color_data = 108'b111010101000111010101000110110010111111111001010101001100100111111011011111111001010101101110100101001010011;
		12'b011000100000: color_data = 108'b110110010111111010101000110101110110111111001010101001010011111111001010111111001010101001100100101000110011;
		12'b011000100001: color_data = 108'b110101110110110110010111111011011101111111001010101000110011111111001010110011001011101001010011111011001100;
		12'b011000100010: color_data = 108'b111011011101110101110110111111111111110011001011111011001100111111001010101111001100101000110011111111111111;
		12'b011000100011: color_data = 108'b111111111111111011011101111111111111101111001100111111111111110011001011101110111011111011001100111111111111;
		12'b011000100100: color_data = 108'b111111111111111111111111111111111111101110111011111111111111101111001100110011001100111111111111111111111111;
		12'b011000100101: color_data = 108'b111111111111111111111111111111111111110011001100111111111111101110111011111011101110111111111111111111111111;
		12'b011000100110: color_data = 108'b111111111111111111111111111111111111111011101110111111111111110011001100111111111111111111111111111111111111;
		12'b011000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111;
		12'b011000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001000101: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111110011001111;
		12'b011001000110: color_data = 108'b111011101111111111111111110011011111111111111111110011001111111111111111111011101111111111111111010001011111;
		12'b011001000111: color_data = 108'b110011011111111011101111010101101110111011101111010001011111111111111111010101101111110011001111001000111011;
		12'b011001001000: color_data = 108'b010101101110110011011111000100111100010101101111001000111011111011101111001000111110010001011111000100101001;
		12'b011001001001: color_data = 108'b000100111100010101101110000100101000001000111110000100101001010101101111001000111100001000111011000100101001;
		12'b011001001010: color_data = 108'b000100101000000100111100000100101001001000111100000100101001001000111110001000111100000100101001000100101001;
		12'b011001001011: color_data = 108'b000100101001000100101000000100101001001000111100000100101001001000111100000100101010000100101001000100101001;
		12'b011001001100: color_data = 108'b000100101001000100101001000100101001000100101010000100101001001000111100000100101000000100101001000100101001;
		12'b011001001101: color_data = 108'b000100101001000100101001000100101001000100101000000100101001000100101010000100101001000100101001000100101001;
		12'b011001001110: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101000000100101001000100101001000100101001;
		12'b011001001111: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b011001010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001;
		12'b011001010001: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101000;
		12'b011001010010: color_data = 108'b000100101001000100101001000100101000000100101001000100101000000100101001000100101001000100101001001000100100;
		12'b011001010011: color_data = 108'b000100101000000100101001000100101000000100101001001000100100000100101001010001000111000100101000000100100110;
		12'b011001010100: color_data = 108'b000100101000000100101000001100111000010001000111000100100110000100101001100001100111001000100100000100101001;
		12'b011001010101: color_data = 108'b001100111000000100101000100101110110100001100111000100101001010001000111110110101000000100100110001000111000;
		12'b011001010110: color_data = 108'b100101110110001100111000110110101000110110101000001000111000100001100111111110111001000100101001100101110110;
		12'b011001010111: color_data = 108'b110110101000100101110110111110111001111110111001100101110110110110101000111111001010001000111000101110000101;
		12'b011001011000: color_data = 108'b111110111001110110101000111110111001111111001010101110000101111110111001111111001010100101110110101110000101;
		12'b011001011001: color_data = 108'b111110111001111110111001111110111001111111001010101110000101111111001010111111001010101110000101101110000101;
		12'b011001011010: color_data = 108'b111110111001111110111001111110111001111111001010101110000101111111001010111111001010101110000101101110000101;
		12'b011001011011: color_data = 108'b111110111001111110111001111110111001111111001010101110000101111111001010111111001010101110000101101110000101;
		12'b011001011100: color_data = 108'b111110111001111110111001111010101000111111001010101110000101111111001010111111001001101110000101101101110101;
		12'b011001011101: color_data = 108'b111010101000111110111001101101110100111111001001101101110101111111001010111010101000101110000101100100010001;
		12'b011001011110: color_data = 108'b101101110100111010101000101001100100111010101000100100010001111111001001111010101000101101110101100100000000;
		12'b011001011111: color_data = 108'b101001100100101101110100101001010011111010101000100100000000111010101000110110010111100100010001101001000100;
		12'b011001100000: color_data = 108'b101001010011101001100100101000110011110110010111101001000100111010101000110101110110100100000000111011011101;
		12'b011001100001: color_data = 108'b101000110011101001010011111011001100110101110110111011011101110110010111111011011101101001000100111111101110;
		12'b011001100010: color_data = 108'b111011001100101000110011111111111111111011011101111111101110110101110110111111111111111011011101111111111111;
		12'b011001100011: color_data = 108'b111111111111111011001100111111111111111111111111111111111111111011011101111111111111111111101110111111111111;
		12'b011001100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010000101: color_data = 108'b111111111111111111111111110011001111111111111111111111111111111111111111111011101111111111111111111011101111;
		12'b011010000110: color_data = 108'b110011001111111111111111010001011111111011101111111011101111111111111111110011011111111111111111101110111111;
		12'b011010000111: color_data = 108'b010001011111110011001111001000111011110011011111101110111111111011101111010101101110111011101111101010111101;
		12'b011010001000: color_data = 108'b001000111011010001011111000100101001010101101110101010111101110011011111000100111100101110111111101010111101;
		12'b011010001001: color_data = 108'b000100101001001000111011000100101001000100111100101010111101010101101110000100101000101010111101101010111101;
		12'b011010001010: color_data = 108'b000100101001000100101001000100101001000100101000101010111101000100111100000100101001101010111101101010111101;
		12'b011010001011: color_data = 108'b000100101001000100101001000100101001000100101001101010111101000100101000000100101001101010111101101110111101;
		12'b011010001100: color_data = 108'b000100101001000100101001000100101001000100101001101110111101000100101001000100101001101010111101011101111011;
		12'b011010001101: color_data = 108'b000100101001000100101001000100101001000100101001011101111011000100101001000100101001101110111101000100101000;
		12'b011010001110: color_data = 108'b000100101001000100101001000100101001000100101001000100101000000100101001000100101001011101111011000100101000;
		12'b011010001111: color_data = 108'b000100101001000100101001000100101001000100101001000100101000000100101001000100101001000100101000000100101001;
		12'b011010010000: color_data = 108'b000100101001000100101001000100101001000100101001000100101001000100101001000100101001000100101000000100101001;
		12'b011010010001: color_data = 108'b000100101001000100101001000100101000000100101001000100101001000100101001000100101001000100101001000100101000;
		12'b011010010010: color_data = 108'b000100101000000100101001001000100100000100101001000100101000000100101001000100101000000100101001000100100111;
		12'b011010010011: color_data = 108'b001000100100000100101000000100100110000100101000000100100111000100101001000100101000000100101000000100100101;
		12'b011010010100: color_data = 108'b000100100110001000100100000100101001000100101000000100100101000100101000001100111000000100100111000100100100;
		12'b011010010101: color_data = 108'b000100101001000100100110001000111000001100111000000100100100000100101000100101110110000100100101000100100100;
		12'b011010010110: color_data = 108'b001000111000000100101001100101110110100101110110000100100100001100111000110110101000000100100100001100110110;
		12'b011010010111: color_data = 108'b100101110110001000111000101110000101110110101000001100110110100101110110111110111001000100100100010001000111;
		12'b011010011000: color_data = 108'b101110000101100101110110101110000101111110111001010001000111110110101000111110111001001100110110010001001000;
		12'b011010011001: color_data = 108'b101110000101101110000101101110000101111110111001010001001000111110111001111110111001010001000111010101011100;
		12'b011010011010: color_data = 108'b101110000101101110000101101110000101111110111001010101011100111110111001111110111001010001001000100000110100;
		12'b011010011011: color_data = 108'b101110000101101110000101101110000101111110111001100000110100111110111001111110111001010101011100100100100001;
		12'b011010011100: color_data = 108'b101110000101101110000101101101110101111110111001100100100001111110111001111010101000100000110100100100100001;
		12'b011010011101: color_data = 108'b101101110101101110000101100100010001111010101000100100100001111110111001101101110100100100100001100000000000;
		12'b011010011110: color_data = 108'b100100010001101101110101100100000000101101110100100000000000111010101000101001100100100100100001101101100110;
		12'b011010011111: color_data = 108'b100100000000100100010001101001000100101001100100101101100110101101110100101001010011100000000000110111001100;
		12'b011010100000: color_data = 108'b101001000100100100000000111011011101101001010011110111001100101001100100101000110011101101100110111111111111;
		12'b011010100001: color_data = 108'b111011011101101001000100111111101110101000110011111111111111101001010011111011001100110111001100111111111111;
		12'b011010100010: color_data = 108'b111111101110111011011101111111111111111011001100111111111111101000110011111111111111111111111111111111111111;
		12'b011010100011: color_data = 108'b111111111111111111101110111111111111111111111111111111111111111011001100111111111111111111111111111111111111;
		12'b011010100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011000101: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111110011001111111111111111111111111111;
		12'b011011000110: color_data = 108'b111011101111111111111111101110111111110011001111111111111111111111111111010001011111111111111111111111111111;
		12'b011011000111: color_data = 108'b101110111111111011101111101010111101010001011111111111111111110011001111001000111011111111111111111111111111;
		12'b011011001000: color_data = 108'b101010111101101110111111101010111101001000111011111111111111010001011111000100101001111111111111111111111111;
		12'b011011001001: color_data = 108'b101010111101101010111101101010111101000100101001111111111111001000111011000100101001111111111111111111111111;
		12'b011011001010: color_data = 108'b101010111101101010111101101010111101000100101001111111111111000100101001000100101001111111111111111111111111;
		12'b011011001011: color_data = 108'b101010111101101010111101101110111101000100101001111111111111000100101001000100101001111111111111111111111111;
		12'b011011001100: color_data = 108'b101110111101101010111101011101111011000100101001111111111111000100101001000100101001111111111111110011001101;
		12'b011011001101: color_data = 108'b011101111011101110111101000100101000000100101001110011001101000100101001000100101001111111111111011001111011;
		12'b011011001110: color_data = 108'b000100101000011101111011000100101000000100101001011001111011000100101001000100101001110011001101011001111011;
		12'b011011001111: color_data = 108'b000100101000000100101000000100101001000100101001011001111011000100101001000100101001011001111011001101001001;
		12'b011011010000: color_data = 108'b000100101001000100101000000100101001000100101001001101001001000100101001000100101001011001111011000100101001;
		12'b011011010001: color_data = 108'b000100101001000100101001000100101000000100101001000100101001000100101001000100101000001101001001000100101001;
		12'b011011010010: color_data = 108'b000100101000000100101001000100100111000100101000000100101001000100101001001000100100000100101001010101011001;
		12'b011011010011: color_data = 108'b000100100111000100101000000100100101001000100100010101011001000100101000000100100110000100101001011101100111;
		12'b011011010100: color_data = 108'b000100100101000100100111000100100100000100100110011101100111001000100100000100101001010101011001011101010101;
		12'b011011010101: color_data = 108'b000100100100000100100101000100100100000100101001011101010101000100100110001000111000011101100111011101010101;
		12'b011011010110: color_data = 108'b000100100100000100100100001100110110001000111000011101010101000100101001100101110110011101010101011001101000;
		12'b011011010111: color_data = 108'b001100110110000100100100010001000111100101110110011001101000001000111000101110000101011101010101010001001010;
		12'b011011011000: color_data = 108'b010001000111001100110110010001001000101110000101010001001010100101110110101110000101011001101000001000111011;
		12'b011011011001: color_data = 108'b010001001000010001000111010101011100101110000101001000111011101110000101101110000101010001001010010101011100;
		12'b011011011010: color_data = 108'b010101011100010001001000100000110100101110000101010101011100101110000101101110000101001000111011100101000110;
		12'b011011011011: color_data = 108'b100000110100010101011100100100100001101110000101100101000110101110000101101110000101010101011100101101000011;
		12'b011011011100: color_data = 108'b100100100001100000110100100100100001101110000101101101000011101110000101101101110101100101000110101101000011;
		12'b011011011101: color_data = 108'b100100100001100100100001100000000000101101110101101101000011101110000101100100010001101101000011100100110010;
		12'b011011011110: color_data = 108'b100000000000100100100001101101100110100100010001100100110010101101110101100100000000101101000011101101110110;
		12'b011011011111: color_data = 108'b101101100110100000000000110111001100100100000000101101110110100100010001101001000100100100110010110110111011;
		12'b011011100000: color_data = 108'b110111001100101101100110111111111111101001000100110110111011100100000000111011011101101101110110111111111111;
		12'b011011100001: color_data = 108'b111111111111110111001100111111111111111011011101111111111111101001000100111111101110110110111011111111111111;
		12'b011011100010: color_data = 108'b111111111111111111111111111111111111111111101110111111111111111011011101111111111111111111111111111111111111;
		12'b011011100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111101110111111111111111111111111111111111111;
		12'b011011100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111;
		12'b011100000110: color_data = 108'b111111111111111111111111111111111111111011101111111111111111111111111111101110111111111111111111111111111111;
		12'b011100000111: color_data = 108'b111111111111111111111111111111111111101110111111111111111111111011101111101010111101111111111111111111111111;
		12'b011100001000: color_data = 108'b111111111111111111111111111111111111101010111101111111111111101110111111101010111101111111111111111111111111;
		12'b011100001001: color_data = 108'b111111111111111111111111111111111111101010111101111111111111101010111101101010111101111111111111111111111111;
		12'b011100001010: color_data = 108'b111111111111111111111111111111111111101010111101111111111111101010111101101010111101111111111111111111111111;
		12'b011100001011: color_data = 108'b111111111111111111111111111111111111101010111101111111111111101010111101101110111101111111111111111111111111;
		12'b011100001100: color_data = 108'b111111111111111111111111110011001101101110111101111111111111101010111101011101111011111111111111111111111111;
		12'b011100001101: color_data = 108'b110011001101111111111111011001111011011101111011111111111111101110111101000100101000111111111111111011101111;
		12'b011100001110: color_data = 108'b011001111011110011001101011001111011000100101000111011101111011101111011000100101000111111111111110111011110;
		12'b011100001111: color_data = 108'b011001111011011001111011001101001001000100101000110111011110000100101000000100101001111011101111011101111011;
		12'b011100010000: color_data = 108'b001101001001011001111011000100101001000100101001011101111011000100101000000100101001110111011110001000111001;
		12'b011100010001: color_data = 108'b000100101001001101001001000100101001000100101001001000111001000100101001000100101000011101111011001101001001;
		12'b011100010010: color_data = 108'b000100101001000100101001010101011001000100101000001101001001000100101001000100100111001000111001110110101001;
		12'b011100010011: color_data = 108'b010101011001000100101001011101100111000100100111110110101001000100101000000100100101001101001001111110111001;
		12'b011100010100: color_data = 108'b011101100111010101011001011101010101000100100101111110111001000100100111000100100100110110101001111110111001;
		12'b011100010101: color_data = 108'b011101010101011101100111011101010101000100100100111110111001000100100101000100100100111110111001111110111001;
		12'b011100010110: color_data = 108'b011101010101011101010101011001101000000100100100111110111001000100100100001100110110111110111001111010111010;
		12'b011100010111: color_data = 108'b011001101000011101010101010001001010001100110110111010111010000100100100010001000111111110111001100110001100;
		12'b011100011000: color_data = 108'b010001001010011001101000001000111011010001000111100110001100001100110110010001001000111010111010010001011101;
		12'b011100011001: color_data = 108'b001000111011010001001010010101011100010001001000010001011101010001000111010101011100100110001100101110000110;
		12'b011100011010: color_data = 108'b010101011100001000111011100101000110010101011100101110000110010001001000100000110100010001011101111010111000;
		12'b011100011011: color_data = 108'b100101000110010101011100101101000011100000110100111010111000010101011100100100100001101110000110111111001010;
		12'b011100011100: color_data = 108'b101101000011100101000110101101000011100100100001111111001010100000110100100100100001111010111000111110111001;
		12'b011100011101: color_data = 108'b101101000011101101000011100100110010100100100001111110111001100100100001100000000000111111001010110010000110;
		12'b011100011110: color_data = 108'b100100110010101101000011101101110110100000000000110010000110100100100001101101100110111110111001101000110010;
		12'b011100011111: color_data = 108'b101101110110100100110010110110111011101101100110101000110010100000000000110111001100110010000110101101010100;
		12'b011100100000: color_data = 108'b110110111011101101110110111111111111110111001100101101010100101101100110111111111111101000110010111111101110;
		12'b011100100001: color_data = 108'b111111111111110110111011111111111111111111111111111111101110110111001100111111111111101101010100111111111111;
		12'b011100100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111111;
		12'b011100100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111110011001101111111111111111111111111;
		12'b011101001101: color_data = 108'b111111111111111111111111111011101111110011001101111111111111111111111111011001111011111111111111110111011110;
		12'b011101001110: color_data = 108'b111011101111111111111111110111011110011001111011110111011110110011001101011001111011111111111111010001011010;
		12'b011101001111: color_data = 108'b110111011110111011101111011101111011011001111011010001011010011001111011001101001001110111011110100110001010;
		12'b011101010000: color_data = 108'b011101111011110111011110001000111001001101001001100110001010011001111011000100101001010001011010111010111001;
		12'b011101010001: color_data = 108'b001000111001011101111011001101001001000100101001111010111001001101001001000100101001100110001010110110101001;
		12'b011101010010: color_data = 108'b001101001001001000111001110110101001000100101001110110101001000100101001010101011001111010111001110010010110;
		12'b011101010011: color_data = 108'b110110101001001101001001111110111001010101011001110010010110000100101001011101100111110110101001110010000101;
		12'b011101010100: color_data = 108'b111110111001110110101001111110111001011101100111110010000101010101011001011101010101110010010110110010000101;
		12'b011101010101: color_data = 108'b111110111001111110111001111110111001011101010101110010000101011101100111011101010101110010000101101110000110;
		12'b011101010110: color_data = 108'b111110111001111110111001111010111010011101010101101110000110011101010101011001101000110010000101011001101101;
		12'b011101010111: color_data = 108'b111010111010111110111001100110001100011001101000011001101101011101010101010001001010101110000110011001101011;
		12'b011101011000: color_data = 108'b100110001100111010111010010001011101010001001010011001101011011001101000001000111011011001101101101110000111;
		12'b011101011001: color_data = 108'b010001011101100110001100101110000110001000111011101110000111010001001010010101011100011001101011111010111001;
		12'b011101011010: color_data = 108'b101110000110010001011101111010111000010101011100111010111001001000111011100101000110101110000111111111001001;
		12'b011101011011: color_data = 108'b111010111000101110000110111111001010100101000110111111001001010101011100101101000011111010111001111111001010;
		12'b011101011100: color_data = 108'b111111001010111010111000111110111001101101000011111111001010100101000110101101000011111111001001111111001010;
		12'b011101011101: color_data = 108'b111110111001111111001010110010000110101101000011111111001010101101000011100100110010111111001010111110111001;
		12'b011101011110: color_data = 108'b110010000110111110111001101000110010100100110010111110111001101101000011101101110110111111001010110010000110;
		12'b011101011111: color_data = 108'b101000110010110010000110101101010100101101110110110010000110100100110010110110111011111110111001110010010111;
		12'b011101100000: color_data = 108'b101101010100101000110010111111101110110110111011110010010111101101110110111111111111110010000110111111111111;
		12'b011101100001: color_data = 108'b111111101110101101010100111111111111111111111111111111111111110110111011111111111111110010010111111111111111;
		12'b011101100010: color_data = 108'b111111111111111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111001101;
		12'b011110001101: color_data = 108'b111111111111111111111111110111011110111111111111101111001101111111111111111011101111111111111111011101111011;
		12'b011110001110: color_data = 108'b110111011110111111111111010001011010111011101111011101111011111111111111110111011110101111001101100110001001;
		12'b011110001111: color_data = 108'b010001011010110111011110100110001010110111011110100110001001111011101111011101111011011101111011110010011000;
		12'b011110010000: color_data = 108'b100110001010010001011010111010111001011101111011110010011000110111011110001000111001100110001001110110010111;
		12'b011110010001: color_data = 108'b111010111001100110001010110110101001001000111001110110010111011101111011001101001001110010011000110010010111;
		12'b011110010010: color_data = 108'b110110101001111010111001110010010110001101001001110010010111001000111001110110101001110110010111011001010111;
		12'b011110010011: color_data = 108'b110010010110110110101001110010000101110110101001011001010111001101001001111110111001110010010111010101000111;
		12'b011110010100: color_data = 108'b110010000101110010010110110010000101111110111001010101000111110110101001111110111001011001010111010101000111;
		12'b011110010101: color_data = 108'b110010000101110010000101101110000110111110111001010101000111111110111001111110111001010101000111010101000111;
		12'b011110010110: color_data = 108'b101110000110110010000101011001101101111110111001010101000111111110111001111010111010010101000111001101001110;
		12'b011110010111: color_data = 108'b011001101101101110000110011001101011111010111010001101001110111110111001100110001100010101000111011001011011;
		12'b011110011000: color_data = 108'b011001101011011001101101101110000111100110001100011001011011111010111010010001011101001101001110110010000101;
		12'b011110011001: color_data = 108'b101110000111011001101011111010111001010001011101110010000101100110001100101110000110011001011011111111001001;
		12'b011110011010: color_data = 108'b111010111001101110000111111111001001101110000110111111001001010001011101111010111000110010000101111111001010;
		12'b011110011011: color_data = 108'b111111001001111010111001111111001010111010111000111111001010101110000110111111001010111111001001111111001010;
		12'b011110011100: color_data = 108'b111111001010111111001001111111001010111111001010111111001010111010111000111110111001111111001010111111001010;
		12'b011110011101: color_data = 108'b111111001010111111001010111110111001111110111001111111001010111111001010110010000110111111001010111111001010;
		12'b011110011110: color_data = 108'b111110111001111111001010110010000110110010000110111111001010111110111001101000110010111111001010110110010111;
		12'b011110011111: color_data = 108'b110010000110111110111001110010010111101000110010110110010111110010000110101101010100111111001010110010101000;
		12'b011110100000: color_data = 108'b110010010111110010000110111111111111101101010100110010101000101000110010111111101110110110010111111111111111;
		12'b011110100001: color_data = 108'b111111111111110010010111111111111111111111101110111111111111101101010100111111111111110010101000111111111111;
		12'b011110100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111101110111111111111111111111111111111111111;
		12'b011110100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b011111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111001100: color_data = 108'b111111111111111111111111101111001101111111111111111111111111111111111111111111111111111111111111100110101100;
		12'b011111001101: color_data = 108'b101111001101111111111111011101111011111111111111100110101100111111111111110111011110111111111111001100111001;
		12'b011111001110: color_data = 108'b011101111011101111001101100110001001110111011110001100111001111111111111010001011010100110101100111010111001;
		12'b011111001111: color_data = 108'b100110001001011101111011110010011000010001011010111010111001110111011110100110001010001100111001110110010110;
		12'b011111010000: color_data = 108'b110010011000100110001001110110010111100110001010110110010110010001011010111010111001111010111001101001110101;
		12'b011111010001: color_data = 108'b110110010111110010011000110010010111111010111001101001110101100110001010110110101001110110010110011101100110;
		12'b011111010010: color_data = 108'b110010010111110110010111011001010111110110101001011101100110111010111001110010010110101001110101001000111000;
		12'b011111010011: color_data = 108'b011001010111110010010111010101000111110010010110001000111000110110101001110010000101011101100110000100101001;
		12'b011111010100: color_data = 108'b010101000111011001010111010101000111110010000101000100101001110010010110110010000101001000111000000100101001;
		12'b011111010101: color_data = 108'b010101000111010101000111010101000111110010000101000100101001110010000101101110000110000100101001000100101001;
		12'b011111010110: color_data = 108'b010101000111010101000111001101001110101110000110000100101001110010000101011001101101000100101001001000111110;
		12'b011111010111: color_data = 108'b001101001110010101000111011001011011011001101101001000111110101110000110011001101011000100101001011001101011;
		12'b011111011000: color_data = 108'b011001011011001101001110110010000101011001101011011001101011011001101101101110000111001000111110110010000101;
		12'b011111011001: color_data = 108'b110010000101011001011011111111001001101110000111110010000101011001101011111010111001011001101011111010101000;
		12'b011111011010: color_data = 108'b111111001001110010000101111111001010111010111001111010101000101110000111111111001001110010000101111110111001;
		12'b011111011011: color_data = 108'b111111001010111111001001111111001010111111001001111110111001111010111001111111001010111010101000111111001010;
		12'b011111011100: color_data = 108'b111111001010111111001010111111001010111111001010111111001010111111001001111111001010111110111001111111001001;
		12'b011111011101: color_data = 108'b111111001010111111001010111111001010111111001010111111001001111111001010111110111001111111001010111010111000;
		12'b011111011110: color_data = 108'b111111001010111111001010110110010111111110111001111010111000111111001010110010000110111111001001110001110101;
		12'b011111011111: color_data = 108'b110110010111111111001010110010101000110010000110110001110101111110111001110010010111111010111000110010000111;
		12'b011111100000: color_data = 108'b110010101000110110010111111111111111110010010111110010000111110010000110111111111111110001110101111111111111;
		12'b011111100001: color_data = 108'b111111111111110010101000111111111111111111111111111111111111110010010111111111111111110010000111111111111111;
		12'b011111100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b011111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b100000001100: color_data = 108'b111111111111111111111111100110101100111111111111111011101111111111111111101111001101111111111111100110011100;
		12'b100000001101: color_data = 108'b100110101100111111111111001100111001101111001101100110011100111111111111011101111011111011101111001100111001;
		12'b100000001110: color_data = 108'b001100111001100110101100111010111001011101111011001100111001101111001101100110001001100110011100110110101001;
		12'b100000001111: color_data = 108'b111010111001001100111001110110010110100110001001110110101001011101111011110010011000001100111001110110010111;
		12'b100000010000: color_data = 108'b110110010110111010111001101001110101110010011000110110010111100110001001110110010111110110101001100001100110;
		12'b100000010001: color_data = 108'b101001110101110110010110011101100110110110010111100001100110110010011000110010010111110110010111001000111001;
		12'b100000010010: color_data = 108'b011101100110101001110101001000111000110010010111001000111001110110010111011001010111100001100110000100101001;
		12'b100000010011: color_data = 108'b001000111000011101100110000100101001011001010111000100101001110010010111010101000111001000111001001000111001;
		12'b100000010100: color_data = 108'b000100101001001000111000000100101001010101000111001000111001011001010111010101000111000100101001001000111001;
		12'b100000010101: color_data = 108'b000100101001000100101001000100101001010101000111001000111001010101000111010101000111001000111001000100101001;
		12'b100000010110: color_data = 108'b000100101001000100101001001000111110010101000111000100101001010101000111001101001110001000111001001000111110;
		12'b100000010111: color_data = 108'b001000111110000100101001011001101011001101001110001000111110010101000111011001011011000100101001011001011011;
		12'b100000011000: color_data = 108'b011001101011001000111110110010000101011001011011011001011011001101001110110010000101001000111110101101110101;
		12'b100000011001: color_data = 108'b110010000101011001101011111010101000110010000101101101110101011001011011111111001001011001011011101110000101;
		12'b100000011010: color_data = 108'b111010101000110010000101111110111001111111001001101110000101110010000101111111001010101101110101111010101000;
		12'b100000011011: color_data = 108'b111110111001111010101000111111001010111111001010111010101000111111001001111111001010101110000101111111001001;
		12'b100000011100: color_data = 108'b111111001010111110111001111111001001111111001010111111001001111111001010111111001010111010101000111110111001;
		12'b100000011101: color_data = 108'b111111001001111111001010111010111000111111001010111110111001111111001010111111001010111111001001101110000101;
		12'b100000011110: color_data = 108'b111010111000111111001001110001110101111111001010101110000101111111001010110110010111111110111001100100100001;
		12'b100000011111: color_data = 108'b110001110101111010111000110010000111110110010111100100100001111111001010110010101000101110000101101001000100;
		12'b100000100000: color_data = 108'b110010000111110001110101111111111111110010101000101001000100110110010111111111111111100100100001111011101110;
		12'b100000100001: color_data = 108'b111111111111110010000111111111111111111111111111111011101110110010101000111111111111101001000100111111111111;
		12'b100000100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111;
		12'b100000100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001001011: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111011110001011;
		12'b100001001100: color_data = 108'b111011101111111111111111100110011100111111111111011110001011111111111111100110101100111111111111001000111001;
		12'b100001001101: color_data = 108'b100110011100111011101111001100111001100110101100001000111001111111111111001100111001011110001011001000111000;
		12'b100001001110: color_data = 108'b001100111001100110011100110110101001001100111001001000111000100110101100111010111001001000111001101110000110;
		12'b100001001111: color_data = 108'b110110101001001100111001110110010111111010111001101110000110001100111001110110010110001000111000111011001010;
		12'b100001010000: color_data = 108'b110110010111110110101001100001100110110110010110111011001010111010111001101001110101101110000110111011101110;
		12'b100001010001: color_data = 108'b100001100110110110010111001000111001101001110101111011101110110110010110011101100110111011001010110011001110;
		12'b100001010010: color_data = 108'b001000111001100001100110000100101001011101100110110011001110101001110101001000111000111011101110011101111001;
		12'b100001010011: color_data = 108'b000100101001001000111001001000111001001000111000011101111001011101100110000100101001110011001110101010101011;
		12'b100001010100: color_data = 108'b001000111001000100101001001000111001000100101001101010101011001000111000000100101001011101111001101110111101;
		12'b100001010101: color_data = 108'b001000111001001000111001000100101001000100101001101110111101000100101001000100101001101010101011011001101001;
		12'b100001010110: color_data = 108'b000100101001001000111001001000111110000100101001011001101001000100101001001000111110101110111101001101001110;
		12'b100001010111: color_data = 108'b001000111110000100101001011001011011001000111110001101001110000100101001011001101011011001101001001101001111;
		12'b100001011000: color_data = 108'b011001011011001000111110101101110101011001101011001101001111001000111110110010000101001101001110010101011100;
		12'b100001011001: color_data = 108'b101101110101011001011011101110000101110010000101010101011100011001101011111010101000001101001111101101110101;
		12'b100001011010: color_data = 108'b101110000101101101110101111010101000111010101000101101110101110010000101111110111001010101011100110010000101;
		12'b100001011011: color_data = 108'b111010101000101110000101111111001001111110111001110010000101111010101000111111001010101101110101110010000110;
		12'b100001011100: color_data = 108'b111111001001111010101000111110111001111111001010110010000110111110111001111111001001110010000101110001110101;
		12'b100001011101: color_data = 108'b111110111001111111001001101110000101111111001001110001110101111111001010111010111000110010000110100100100001;
		12'b100001011110: color_data = 108'b101110000101111110111001100100100001111010111000100100100001111111001001110001110101110001110101010100010001;
		12'b100001011111: color_data = 108'b100100100001101110000101101001000100110001110101010100010001111010111000110010000111100100100001010000110011;
		12'b100001100000: color_data = 108'b101001000100100100100001111011101110110010000111010000110011110001110101111111111111010100010001011101110111;
		12'b100001100001: color_data = 108'b111011101110101001000100111111111111111111111111011101110111110010000111111111111111010000110011110111011101;
		12'b100001100010: color_data = 108'b111111111111111011101110111111111111111111111111110111011101111111111111111111111111011101110111111111111111;
		12'b100001100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101111111111111;
		12'b100001100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b100010001011: color_data = 108'b111111111111111111111111011110001011111111111111111011101111111111111111111011101111111111111111010101101010;
		12'b100010001100: color_data = 108'b011110001011111111111111001000111001111011101111010101101010111111111111100110011100111011101111000100101000;
		12'b100010001101: color_data = 108'b001000111001011110001011001000111000100110011100000100101000111011101111001100111001010101101010001000101000;
		12'b100010001110: color_data = 108'b001000111000001000111001101110000110001100111001001000101000100110011100110110101001000100101000100100110011;
		12'b100010001111: color_data = 108'b101110000110001000111000111011001010110110101001100100110011001100111001110110010111001000101000111010111011;
		12'b100010010000: color_data = 108'b111011001010101110000110111011101110110110010111111010111011110110101001100001100110100100110011111011111111;
		12'b100010010001: color_data = 108'b111011101110111011001010110011001110100001100110111011111111110110010111001000111001111010111011110011001100;
		12'b100010010010: color_data = 108'b110011001110111011101110011101111001001000111001110011001100100001100110000100101001111011111111110011001100;
		12'b100010010011: color_data = 108'b011101111001110011001110101010101011000100101001110011001100001000111001001000111001110011001100111011101110;
		12'b100010010100: color_data = 108'b101010101011011101111001101110111101001000111001111011101110000100101001001000111001110011001100111111111111;
		12'b100010010101: color_data = 108'b101110111101101010101011011001101001001000111001111111111111001000111001000100101001111011101110101110111100;
		12'b100010010110: color_data = 108'b011001101001101110111101001101001110000100101001101110111100001000111001001000111110111111111111010001011100;
		12'b100010010111: color_data = 108'b001101001110011001101001001101001111001000111110010001011100000100101001011001011011101110111100001000111110;
		12'b100010011000: color_data = 108'b001101001111001101001110010101011100011001011011001000111110001000111110101101110101010001011100001101001111;
		12'b100010011001: color_data = 108'b010101011100001101001111101101110101101101110101001101001111011001011011101110000101001000111110011001101011;
		12'b100010011010: color_data = 108'b101101110101010101011100110010000101101110000101011001101011101101110101111010101000001101001111011001101010;
		12'b100010011011: color_data = 108'b110010000101101101110101110010000110111010101000011001101010101110000101111111001001011001101011011001101010;
		12'b100010011100: color_data = 108'b110010000110110010000101110001110101111111001001011001101010111010101000111110111001011001101010011001011010;
		12'b100010011101: color_data = 108'b110001110101110010000110100100100001111110111001011001011010111111001001101110000101011001101010010100010101;
		12'b100010011110: color_data = 108'b100100100001110001110101010100010001101110000101010100010101111110111001100100100001011001011010010000100100;
		12'b100010011111: color_data = 108'b010100010001100100100001010000110011100100100001010000100100101110000101101001000100010100010101010001000100;
		12'b100010100000: color_data = 108'b010000110011010100010001011101110111101001000100010001000100100100100001111011101110010000100100011001100111;
		12'b100010100001: color_data = 108'b011101110111010000110011110111011101111011101110011001100111101001000100111111111111010001000100101010101011;
		12'b100010100010: color_data = 108'b110111011101011101110111111111111111111111111111101010101011111011101110111111111111011001100111110111011101;
		12'b100010100011: color_data = 108'b111111111111110111011101111111111111111111111111110111011101111111111111111111111111101010101011111111111111;
		12'b100010100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101111111111111;
		12'b100010100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011001010: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b100011001011: color_data = 108'b111011101111111111111111010101101010111111111111111011101111111111111111011110001011111111111111010101101010;
		12'b100011001100: color_data = 108'b010101101010111011101111000100101000011110001011010101101010111111111111001000111001111011101111000100101001;
		12'b100011001101: color_data = 108'b000100101000010101101010001000101000001000111001000100101001011110001011001000111000010101101010001000101000;
		12'b100011001110: color_data = 108'b001000101000000100101000100100110011001000111000001000101000001000111001101110000110000100101001011000000010;
		12'b100011001111: color_data = 108'b100100110011001000101000111010111011101110000110011000000010001000111000111011001010001000101000101110011001;
		12'b100011010000: color_data = 108'b111010111011100100110011111011111111111011001010101110011001101110000110111011101110011000000010110011001100;
		12'b100011010001: color_data = 108'b111011111111111010111011110011001100111011101110110011001100111011001010110011001110101110011001011101111000;
		12'b100011010010: color_data = 108'b110011001100111011111111110011001100110011001110011101111000111011101110011101111001110011001100110011001101;
		12'b100011010011: color_data = 108'b110011001100110011001100111011101110011101111001110011001101110011001110101010101011011101111000111011101110;
		12'b100011010100: color_data = 108'b111011101110110011001100111111111111101010101011111011101110011101111001101110111101110011001101111011101110;
		12'b100011010101: color_data = 108'b111111111111111011101110101110111100101110111101111011101110101010101011011001101001111011101110110111011110;
		12'b100011010110: color_data = 108'b101110111100111111111111010001011100011001101001110111011110101110111101001101001110111011101110010001011010;
		12'b100011010111: color_data = 108'b010001011100101110111100001000111110001101001110010001011010011001101001001101001111110111011110000100111100;
		12'b100011011000: color_data = 108'b001000111110010001011100001101001111001101001111000100111100001101001110010101011100010001011010001001001111;
		12'b100011011001: color_data = 108'b001101001111001000111110011001101011010101011100001001001111001101001111101101110101000100111100001000111110;
		12'b100011011010: color_data = 108'b011001101011001101001111011001101010101101110101001000111110010101011100110010000101001001001111001000111101;
		12'b100011011011: color_data = 108'b011001101010011001101011011001101010110010000101001000111101101101110101110010000110001000111110001000111101;
		12'b100011011100: color_data = 108'b011001101010011001101010011001011010110010000110001000111101110010000101110001110101001000111101001000111101;
		12'b100011011101: color_data = 108'b011001011010011001101010010100010101110001110101001000111101110010000110100100100001001000111101000100101000;
		12'b100011011110: color_data = 108'b010100010101011001011010010000100100100100100001000100101000110001110101010100010001001000111101001100110110;
		12'b100011011111: color_data = 108'b010000100100010100010101010001000100010100010001001100110110100100100001010000110011000100101000010101010110;
		12'b100011100000: color_data = 108'b010001000100010000100100011001100111010000110011010101010110010100010001011101110111001100110110011101111001;
		12'b100011100001: color_data = 108'b011001100111010001000100101010101011011101110111011101111001010000110011110111011101010101010110011101111000;
		12'b100011100010: color_data = 108'b101010101011011001100111110111011101110111011101011101111000011101110111111111111111011101111001101110111100;
		12'b100011100011: color_data = 108'b110111011101101010101011111111111111111111111111101110111100110111011101111111111111011101111000111111111111;
		12'b100011100100: color_data = 108'b111111111111110111011101111111111111111111111111111111111111111111111111111111111111101110111100111111111111;
		12'b100011100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100001010: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111011101111111111111111111011101111;
		12'b100100001011: color_data = 108'b111011101111111111111111010101101010111011101111111011101111111111111111010101101010111111111111010101101010;
		12'b100100001100: color_data = 108'b010101101010111011101111000100101001010101101010010101101010111011101111000100101000111011101111000100101001;
		12'b100100001101: color_data = 108'b000100101001010101101010001000101000000100101000000100101001010101101010001000101000010101101010000100101001;
		12'b100100001110: color_data = 108'b001000101000000100101001011000000010001000101000000100101001000100101000100100110011000100101001001000101000;
		12'b100100001111: color_data = 108'b011000000010001000101000101110011001100100110011001000101000001000101000111010111011000100101001011001101001;
		12'b100100010000: color_data = 108'b101110011001011000000010110011001100111010111011011001101001100100110011111011111111001000101000011101111000;
		12'b100100010001: color_data = 108'b110011001100101110011001011101111000111011111111011101111000111010111011110011001100011001101001010101010110;
		12'b100100010010: color_data = 108'b011101111000110011001100110011001101110011001100010101010110111011111111110011001100011101111000011101111000;
		12'b100100010011: color_data = 108'b110011001101011101111000111011101110110011001100011101111000110011001100111011101110010101010110100010001001;
		12'b100100010100: color_data = 108'b111011101110110011001101111011101110111011101110100010001001110011001100111111111111011101111000100010001001;
		12'b100100010101: color_data = 108'b111011101110111011101110110111011110111111111111100010001001111011101110101110111100100010001001100010001001;
		12'b100100010110: color_data = 108'b110111011110111011101110010001011010101110111100100010001001111111111111010001011100100010001001001100111001;
		12'b100100010111: color_data = 108'b010001011010110111011110000100111100010001011100001100111001101110111100001000111110100010001001000100111100;
		12'b100100011000: color_data = 108'b000100111100010001011010001001001111001000111110000100111100010001011100001101001111001100111001001001001110;
		12'b100100011001: color_data = 108'b001001001111000100111100001000111110001101001111001001001110001000111110011001101011000100111100001000111001;
		12'b100100011010: color_data = 108'b001000111110001001001111001000111101011001101011001000111001001101001111011001101010001001001110001000100101;
		12'b100100011011: color_data = 108'b001000111101001000111110001000111101011001101010001000100101011001101011011001101010001000111001001000100101;
		12'b100100011100: color_data = 108'b001000111101001000111101001000111101011001101010001000100101011001101010011001011010001000100101000100101000;
		12'b100100011101: color_data = 108'b001000111101001000111101000100101000011001011010000100101000011001101010010100010101001000100101001000100011;
		12'b100100011110: color_data = 108'b000100101000001000111101001100110110010100010101001000100011011001011010010000100100000100101000001100110100;
		12'b100100011111: color_data = 108'b001100110110000100101000010101010110010000100100001100110100010100010101010001000100001000100011010101010110;
		12'b100100100000: color_data = 108'b010101010110001100110110011101111001010001000100010101010110010000100100011001100111001100110100011101111000;
		12'b100100100001: color_data = 108'b011101111001010101010110011101111000011001100111011101111000010001000100101010101011010101010110100010001001;
		12'b100100100010: color_data = 108'b011101111000011101111001101110111100101010101011100010001001011001100111110111011101011101111000101110111100;
		12'b100100100011: color_data = 108'b101110111100011101111000111111111111110111011101101110111100101010101011111111111111100010001001111111111111;
		12'b100100100100: color_data = 108'b111111111111101110111100111111111111111111111111111111111111110111011101111111111111101110111100111111111111;
		12'b100100100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101001010: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111011101111111111111111111011101111;
		12'b100101001011: color_data = 108'b111011101111111111111111010101101010111011101111111011101111111111111111010101101010111111111111010101101010;
		12'b100101001100: color_data = 108'b010101101010111011101111000100101001010101101010010101101010111011101111000100101001111011101111010001011010;
		12'b100101001101: color_data = 108'b000100101001010101101010000100101001000100101001010001011010010101101010001000101000010101101010101110111101;
		12'b100101001110: color_data = 108'b000100101001000100101001001000101000001000101000101110111101000100101001011000000010010001011010101110111101;
		12'b100101001111: color_data = 108'b001000101000000100101001011001101001011000000010101110111101001000101000101110011001101110111101110011001101;
		12'b100101010000: color_data = 108'b011001101001001000101000011101111000101110011001110011001101011000000010110011001100101110111101101110111011;
		12'b100101010001: color_data = 108'b011101111000011001101001010101010110110011001100101110111011101110011001011101111000110011001101011101111000;
		12'b100101010010: color_data = 108'b010101010110011101111000011101111000011101111000011101111000110011001100110011001101101110111011011101111000;
		12'b100101010011: color_data = 108'b011101111000010101010110100010001001110011001101011101111000011101111000111011101110011101111000011101111001;
		12'b100101010100: color_data = 108'b100010001001011101111000100010001001111011101110011101111001110011001101111011101110011101111000011101111001;
		12'b100101010101: color_data = 108'b100010001001100010001001100010001001111011101110011101111001111011101110110111011110011101111001011101111001;
		12'b100101010110: color_data = 108'b100010001001100010001001001100111001110111011110011101111001111011101110010001011010011101111001010101101100;
		12'b100101010111: color_data = 108'b001100111001100010001001000100111100010001011010010101101100110111011110000100111100011101111001001101011111;
		12'b100101011000: color_data = 108'b000100111100001100111001001001001110000100111100001101011111010001011010001001001111010101101100010001011111;
		12'b100101011001: color_data = 108'b001001001110000100111100001000111001001001001111010001011111000100111100001000111110001101011111101010111101;
		12'b100101011010: color_data = 108'b001000111001001001001110001000100101001000111110101010111101001001001111001000111101010001011111010001011001;
		12'b100101011011: color_data = 108'b001000100101001000111001001000100101001000111101010001011001001000111110001000111101101010111101000100100111;
		12'b100101011100: color_data = 108'b001000100101001000100101000100101000001000111101000100100111001000111101001000111101010001011001000100101000;
		12'b100101011101: color_data = 108'b000100101000001000100101001000100011001000111101000100101000001000111101000100101000000100100111001000100010;
		12'b100101011110: color_data = 108'b001000100011000100101000001100110100000100101000001000100010001000111101001100110110000100101000001000100010;
		12'b100101011111: color_data = 108'b001100110100001000100011010101010110001100110110001000100010000100101000010101010110001000100010001100110011;
		12'b100101100000: color_data = 108'b010101010110001100110100011101111000010101010110001100110011001100110110011101111001001000100010010101010110;
		12'b100101100001: color_data = 108'b011101111000010101010110100010001001011101111001010101010110010101010110011101111000001100110011101110111100;
		12'b100101100010: color_data = 108'b100010001001011101111000101110111100011101111000101110111100011101111001101110111100010101010110111011101110;
		12'b100101100011: color_data = 108'b101110111100100010001001111111111111101110111100111011101110011101111000111111111111101110111100111111111111;
		12'b100101100100: color_data = 108'b111111111111101110111100111111111111111111111111111111111111101110111100111111111111111011101110111111111111;
		12'b100101100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110001010: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111011101111111111111111111111111111;
		12'b100110001011: color_data = 108'b111011101111111111111111010101101010111011101111111111111111111111111111010101101010111111111111100110011100;
		12'b100110001100: color_data = 108'b010101101010111011101111010001011010010101101010100110011100111011101111000100101001111111111111101010101101;
		12'b100110001101: color_data = 108'b010001011010010101101010101110111101000100101001101010101101010101101010000100101001100110011100111111111111;
		12'b100110001110: color_data = 108'b101110111101010001011010101110111101000100101001111111111111000100101001001000101000101010101101111111111111;
		12'b100110001111: color_data = 108'b101110111101101110111101110011001101001000101000111111111111000100101001011001101001111111111111111111111111;
		12'b100110010000: color_data = 108'b110011001101101110111101101110111011011001101001111111111111001000101000011101111000111111111111111011011110;
		12'b100110010001: color_data = 108'b101110111011110011001101011101111000011101111000111011011110011001101001010101010110111111111111101010101011;
		12'b100110010010: color_data = 108'b011101111000101110111011011101111000010101010110101010101011011101111000011101111000111011011110100010001001;
		12'b100110010011: color_data = 108'b011101111000011101111000011101111001011101111000100010001001010101010110100010001001101010101011011101111000;
		12'b100110010100: color_data = 108'b011101111001011101111000011101111001100010001001011101111000011101111000100010001001100010001001011101111000;
		12'b100110010101: color_data = 108'b011101111001011101111001011101111001100010001001011101111000100010001001100010001001011101111000010101011001;
		12'b100110010110: color_data = 108'b011101111001011101111001010101101100100010001001010101011001100010001001001100111001011101111000010101111110;
		12'b100110010111: color_data = 108'b010101101100011101111001001101011111001100111001010101111110100010001001000100111100010101011001011110001111;
		12'b100110011000: color_data = 108'b001101011111010101101100010001011111000100111100011110001111001100111001001001001110010101111110100110101111;
		12'b100110011001: color_data = 108'b010001011111001101011111101010111101001001001110100110101111000100111100001000111001011110001111111011101111;
		12'b100110011010: color_data = 108'b101010111101010001011111010001011001001000111001111011101111001001001110001000100101100110101111010101101011;
		12'b100110011011: color_data = 108'b010001011001101010111101000100100111001000100101010101101011001000111001001000100101111011101111000100101001;
		12'b100110011100: color_data = 108'b000100100111010001011001000100101000001000100101000100101001001000100101000100101000010101101011001000111000;
		12'b100110011101: color_data = 108'b000100101000000100100111001000100010000100101000001000111000001000100101001000100011000100101001011101110111;
		12'b100110011110: color_data = 108'b001000100010000100101000001000100010001000100011011101110111000100101000001100110100001000111000011101110111;
		12'b100110011111: color_data = 108'b001000100010001000100010001100110011001100110100011101110111001000100011010101010110011101110111100010001000;
		12'b100110100000: color_data = 108'b001100110011001000100010010101010110010101010110100010001000001100110100011101111000011101110111100110011001;
		12'b100110100001: color_data = 108'b010101010110001100110011101110111100011101111000100110011001010101010110100010001001100010001000111011101110;
		12'b100110100010: color_data = 108'b101110111100010101010110111011101110100010001001111011101110011101111000101110111100100110011001111111111111;
		12'b100110100011: color_data = 108'b111011101110101110111100111111111111101110111100111111111111100010001001111111111111111011101110111111111111;
		12'b100110100100: color_data = 108'b111111111111111011101110111111111111111111111111111111111111101110111100111111111111111111111111111111111111;
		12'b100110100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b100111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111111111111111;
		12'b100111001011: color_data = 108'b111111111111111111111111100110011100111011101111111111111111111111111111010101101010111111111111111111111111;
		12'b100111001100: color_data = 108'b100110011100111111111111101010101101010101101010111111111111111011101111010001011010111111111111111111111111;
		12'b100111001101: color_data = 108'b101010101101100110011100111111111111010001011010111111111111010101101010101110111101111111111111111111111111;
		12'b100111001110: color_data = 108'b111111111111101010101101111111111111101110111101111111111111010001011010101110111101111111111111111111111111;
		12'b100111001111: color_data = 108'b111111111111111111111111111111111111101110111101111111111111101110111101110011001101111111111111111111111111;
		12'b100111010000: color_data = 108'b111111111111111111111111111011011110110011001101111111111111101110111101101110111011111111111111111111111111;
		12'b100111010001: color_data = 108'b111011011110111111111111101010101011101110111011111111111111110011001101011101111000111111111111111011101110;
		12'b100111010010: color_data = 108'b101010101011111011011110100010001001011101111000111011101110101110111011011101111000111111111111101010101010;
		12'b100111010011: color_data = 108'b100010001001101010101011011101111000011101111000101010101010011101111000011101111001111011101110100110011001;
		12'b100111010100: color_data = 108'b011101111000100010001001011101111000011101111001100110011001011101111000011101111001101010101010011101111001;
		12'b100111010101: color_data = 108'b011101111000011101111000010101011001011101111001011101111001011101111001011101111001100110011001000100101001;
		12'b100111010110: color_data = 108'b010101011001011101111000010101111110011101111001000100101001011101111001010101101100011101111001010001101110;
		12'b100111010111: color_data = 108'b010101111110010101011001011110001111010101101100010001101110011101111001001101011111000100101001101010111111;
		12'b100111011000: color_data = 108'b011110001111010101111110100110101111001101011111101010111111010101101100010001011111010001101110111111111111;
		12'b100111011001: color_data = 108'b100110101111011110001111111011101111010001011111111111111111001101011111101010111101101010111111111011101111;
		12'b100111011010: color_data = 108'b111011101111100110101111010101101011101010111101111011101111010001011111010001011001111111111111010101101010;
		12'b100111011011: color_data = 108'b010101101011111011101111000100101001010001011001010101101010101010111101000100100111111011101111000100101000;
		12'b100111011100: color_data = 108'b000100101001010101101011001000111000000100100111000100101000010001011001000100101000010101101010001101001001;
		12'b100111011101: color_data = 108'b001000111000000100101001011101110111000100101000001101001001000100100111001000100010000100101000110111011110;
		12'b100111011110: color_data = 108'b011101110111001000111000011101110111001000100010110111011110000100101000001000100010001101001001111111111111;
		12'b100111011111: color_data = 108'b011101110111011101110111100010001000001000100010111111111111001000100010001100110011110111011110111111111111;
		12'b100111100000: color_data = 108'b100010001000011101110111100110011001001100110011111111111111001000100010010101010110111111111111111111111111;
		12'b100111100001: color_data = 108'b100110011001100010001000111011101110010101010110111111111111001100110011101110111100111111111111111111111111;
		12'b100111100010: color_data = 108'b111011101110100110011001111111111111101110111100111111111111010101010110111011101110111111111111111111111111;
		12'b100111100011: color_data = 108'b111111111111111011101110111111111111111011101110111111111111101110111100111111111111111111111111111111111111;
		12'b100111100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111;
		12'b100111100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b100111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111100110011100111111111111111111111111;
		12'b101000001100: color_data = 108'b111111111111111111111111111111111111100110011100111111111111111111111111101010101101111111111111111111111111;
		12'b101000001101: color_data = 108'b111111111111111111111111111111111111101010101101111111111111100110011100111111111111111111111111111111111111;
		12'b101000001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111101010101101111111111111111111111111111111111111;
		12'b101000001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000010000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011011110111111111111111111111111;
		12'b101000010001: color_data = 108'b111111111111111111111111111011101110111011011110111111111111111111111111101010101011111111111111111111111111;
		12'b101000010010: color_data = 108'b111011101110111111111111101010101010101010101011111111111111111011011110100010001001111111111111111011101110;
		12'b101000010011: color_data = 108'b101010101010111011101110100110011001100010001001111011101110101010101011011101111000111111111111111011101110;
		12'b101000010100: color_data = 108'b100110011001101010101010011101111001011101111000111011101110100010001001011101111000111011101110101110111101;
		12'b101000010101: color_data = 108'b011101111001100110011001000100101001011101111000101110111101011101111000010101011001111011101110001000111001;
		12'b101000010110: color_data = 108'b000100101001011101111001010001101110010101011001001000111001011101111000010101111110101110111101010001101110;
		12'b101000010111: color_data = 108'b010001101110000100101001101010111111010101111110010001101110010101011001011110001111001000111001101010111111;
		12'b101000011000: color_data = 108'b101010111111010001101110111111111111011110001111101010111111010101111110100110101111010001101110111111111111;
		12'b101000011001: color_data = 108'b111111111111101010111111111011101111100110101111111111111111011110001111111011101111101010111111111011101111;
		12'b101000011010: color_data = 108'b111011101111111111111111010101101010111011101111111011101111100110101111010101101011111111111111010101101010;
		12'b101000011011: color_data = 108'b010101101010111011101111000100101000010101101011010101101010111011101111000100101001111011101111000100101000;
		12'b101000011100: color_data = 108'b000100101000010101101010001101001001000100101001000100101000010101101011001000111000010101101010001101001001;
		12'b101000011101: color_data = 108'b001101001001000100101000110111011110001000111000001101001001000100101001011101110111000100101000110111011110;
		12'b101000011110: color_data = 108'b110111011110001101001001111111111111011101110111110111011110001000111000011101110111001101001001111111111111;
		12'b101000011111: color_data = 108'b111111111111110111011110111111111111011101110111111111111111011101110111100010001000110111011110111111111111;
		12'b101000100000: color_data = 108'b111111111111111111111111111111111111100010001000111111111111011101110111100110011001111111111111111111111111;
		12'b101000100001: color_data = 108'b111111111111111111111111111111111111100110011001111111111111100010001000111011101110111111111111111111111111;
		12'b101000100010: color_data = 108'b111111111111111111111111111111111111111011101110111111111111100110011001111111111111111111111111111111111111;
		12'b101000100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111;
		12'b101000100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001010000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001010001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111;
		12'b101001010010: color_data = 108'b111111111111111111111111111011101110111011101110111111111111111111111111101010101010111111111111111111111111;
		12'b101001010011: color_data = 108'b111011101110111111111111111011101110101010101010111111111111111011101110100110011001111111111111101010101100;
		12'b101001010100: color_data = 108'b111011101110111011101110101110111101100110011001101010101100101010101010011101111001111111111111010101101011;
		12'b101001010101: color_data = 108'b101110111101111011101110001000111001011101111001010101101011100110011001000100101001101010101100010001101101;
		12'b101001010110: color_data = 108'b001000111001101110111101010001101110000100101001010001101101011101111001010001101110010101101011101010111110;
		12'b101001010111: color_data = 108'b010001101110001000111001101010111111010001101110101010111110000100101001101010111111010001101101110111011111;
		12'b101001011000: color_data = 108'b101010111111010001101110111111111111101010111111110111011111010001101110111111111111101010111110111111111111;
		12'b101001011001: color_data = 108'b111111111111101010111111111011101111111111111111111111111111101010111111111011101111110111011111111011101111;
		12'b101001011010: color_data = 108'b111011101111111111111111010101101010111011101111111011101111111111111111010101101010111111111111010101101010;
		12'b101001011011: color_data = 108'b010101101010111011101111000100101000010101101010010101101010111011101111000100101000111011101111000100101000;
		12'b101001011100: color_data = 108'b000100101000010101101010001101001001000100101000000100101000010101101010001101001001010101101010001101001001;
		12'b101001011101: color_data = 108'b001101001001000100101000110111011110001101001001001101001001000100101000110111011110000100101000110111011110;
		12'b101001011110: color_data = 108'b110111011110001101001001111111111111110111011110110111011110001101001001111111111111001101001001111111111111;
		12'b101001011111: color_data = 108'b111111111111110111011110111111111111111111111111111111111111110111011110111111111111110111011110111111111111;
		12'b101001100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010010000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010010001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010010010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111;
		12'b101010010011: color_data = 108'b111111111111111111111111101010101100111011101110111111111111111111111111111011101110111111111111011110001011;
		12'b101010010100: color_data = 108'b101010101100111111111111010101101011111011101110011110001011111011101110101110111101111111111111001000111010;
		12'b101010010101: color_data = 108'b010101101011101010101100010001101101101110111101001000111010111011101110001000111001011110001011011001111111;
		12'b101010010110: color_data = 108'b010001101101010101101011101010111110001000111001011001111111101110111101010001101110001000111010110111011111;
		12'b101010010111: color_data = 108'b101010111110010001101101110111011111010001101110110111011111001000111001101010111111011001111111111111111111;
		12'b101010011000: color_data = 108'b110111011111101010111110111111111111101010111111111111111111010001101110111111111111110111011111111111111111;
		12'b101010011001: color_data = 108'b111111111111110111011111111011101111111111111111111111111111101010111111111011101111111111111111111111111111;
		12'b101010011010: color_data = 108'b111011101111111111111111010101101010111011101111111111111111111111111111010101101010111111111111010101101010;
		12'b101010011011: color_data = 108'b010101101010111011101111000100101000010101101010010101101010111011101111000100101000111111111111000100101000;
		12'b101010011100: color_data = 108'b000100101000010101101010001101001001000100101000000100101000010101101010001101001001010101101010001100111001;
		12'b101010011101: color_data = 108'b001101001001000100101000110111011110001101001001001100111001000100101000110111011110000100101000110111011110;
		12'b101010011110: color_data = 108'b110111011110001101001001111111111111110111011110110111011110001101001001111111111111001100111001111111111111;
		12'b101010011111: color_data = 108'b111111111111110111011110111111111111111111111111111111111111110111011110111111111111110111011110111111111111;
		12'b101010100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011010000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111;
		12'b101011010001: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111111111111111011101110;
		12'b101011010010: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111011101111111011101110;
		12'b101011010011: color_data = 108'b111111111111111111111111011110001011111111111111111011101110111111111111101010101100111011101110100010001100;
		12'b101011010100: color_data = 108'b011110001011111111111111001000111010101010101100100010001100111111111111010101101011111011101110001101001011;
		12'b101011010101: color_data = 108'b001000111010011110001011011001111111010101101011001101001011101010101100010001101101100010001100011110001111;
		12'b101011010110: color_data = 108'b011001111111001000111010110111011111010001101101011110001111010101101011101010111110001101001011110111011111;
		12'b101011010111: color_data = 108'b110111011111011001111111111111111111101010111110110111011111010001101101110111011111011110001111111111111111;
		12'b101011011000: color_data = 108'b111111111111110111011111111111111111110111011111111111111111101010111110111111111111110111011111111011101110;
		12'b101011011001: color_data = 108'b111111111111111111111111111111111111111111111111111011101110110111011111111011101111111111111111111011101110;
		12'b101011011010: color_data = 108'b111111111111111111111111010101101010111011101111111011101110111111111111010101101010111011101110010101101010;
		12'b101011011011: color_data = 108'b010101101010111111111111000100101000010101101010010101101010111011101111000100101000111011101110000100101000;
		12'b101011011100: color_data = 108'b000100101000010101101010001100111001000100101000000100101000010101101010001101001001010101101010001101001001;
		12'b101011011101: color_data = 108'b001100111001000100101000110111011110001101001001001101001001000100101000110111011110000100101000110011011101;
		12'b101011011110: color_data = 108'b110111011110001100111001111111111111110111011110110011011101001101001001111111111111001101001001111111111111;
		12'b101011011111: color_data = 108'b111111111111110111011110111111111111111111111111111111111111110111011110111111111111110011011101111111111111;
		12'b101011100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100010000: color_data = 108'b111111111111111111111111111011101111111111111111111111111111111111111111111111111111111111111111110111011101;
		12'b101100010001: color_data = 108'b111011101111111111111111111011101110111111111111110111011101111111111111111111111111111111111111100110011010;
		12'b101100010010: color_data = 108'b111011101110111011101111111011101110111111111111100110011010111111111111111111111111110111011101101110111100;
		12'b101100010011: color_data = 108'b111011101110111011101110100010001100111111111111101110111100111111111111011110001011100110011010110011001101;
		12'b101100010100: color_data = 108'b100010001100111011101110001101001011011110001011110011001101111111111111001000111010101110111100110111011110;
		12'b101100010101: color_data = 108'b001101001011100010001100011110001111001000111010110111011110011110001011011001111111110011001101110111101111;
		12'b101100010110: color_data = 108'b011110001111001101001011110111011111011001111111110111101111001000111010110111011111110111011110111011101111;
		12'b101100010111: color_data = 108'b110111011111011110001111111111111111110111011111111011101111011001111111111111111111110111101111111111111111;
		12'b101100011000: color_data = 108'b111111111111110111011111111011101110111111111111111111111111110111011111111111111111111011101111110111011101;
		12'b101100011001: color_data = 108'b111011101110111111111111111011101110111111111111110111011101111111111111111111111111111111111111011001100111;
		12'b101100011010: color_data = 108'b111011101110111011101110010101101010111111111111011001100111111111111111010101101010110111011101011001101000;
		12'b101100011011: color_data = 108'b010101101010111011101110000100101000010101101010011001101000111111111111000100101000011001100111011101111001;
		12'b101100011100: color_data = 108'b000100101000010101101010001101001001000100101000011101111001010101101010001100111001011001101000011101111001;
		12'b101100011101: color_data = 108'b001101001001000100101000110011011101001100111001011101111001000100101000110111011110011101111001100010001001;
		12'b101100011110: color_data = 108'b110011011101001101001001111111111111110111011110100010001001001100111001111111111111011101111001110011001101;
		12'b101100011111: color_data = 108'b111111111111110011011101111111111111111111111111110011001101110111011110111111111111100010001001111111111111;
		12'b101100100000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001101111111111111;
		12'b101100100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101010000: color_data = 108'b111111111111111111111111110111011101111111111111111111111111111111111111111011101111111111111111110111011101;
		12'b101101010001: color_data = 108'b110111011101111111111111100110011010111011101111110111011101111111111111111011101110111111111111100010001001;
		12'b101101010010: color_data = 108'b100110011010110111011101101110111100111011101110100010001001111011101111111011101110110111011101100110011010;
		12'b101101010011: color_data = 108'b101110111100100110011010110011001101111011101110100110011010111011101110100010001100100010001001101010101011;
		12'b101101010100: color_data = 108'b110011001101101110111100110111011110100010001100101010101011111011101110001101001011100110011010101110111100;
		12'b101101010101: color_data = 108'b110111011110110011001101110111101111001101001011101110111100100010001100011110001111101010101011110111011110;
		12'b101101010110: color_data = 108'b110111101111110111011110111011101111011110001111110111011110001101001011110111011111101110111100110111011110;
		12'b101101010111: color_data = 108'b111011101111110111101111111111111111110111011111110111011110011110001111111111111111110111011110111011101110;
		12'b101101011000: color_data = 108'b111111111111111011101111110111011101111111111111111011101110110111011111111011101110110111011110110111011101;
		12'b101101011001: color_data = 108'b110111011101111111111111011001100111111011101110110111011101111111111111111011101110111011101110010101010110;
		12'b101101011010: color_data = 108'b011001100111110111011101011001101000111011101110010101010110111011101110010101101010110111011101010101010110;
		12'b101101011011: color_data = 108'b011001101000011001100111011101111001010101101010010101010110111011101110000100101000010101010110011001100110;
		12'b101101011100: color_data = 108'b011101111001011001101000011101111001000100101000011001100110010101101010001101001001010101010110011001100111;
		12'b101101011101: color_data = 108'b011101111001011101111001100010001001001101001001011001100111000100101000110011011101011001100110011101111000;
		12'b101101011110: color_data = 108'b100010001001011101111001110011001101110011011101011101111000001101001001111111111111011001100111100110011010;
		12'b101101011111: color_data = 108'b110011001101100010001001111111111111111111111111100110011010110011011101111111111111011101111000110011001100;
		12'b101101100000: color_data = 108'b111111111111110011001101111111111111111111111111110011001100111111111111111111111111100110011010111111111111;
		12'b101101100001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001100111111111111;
		12'b101101100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110001111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101;
		12'b101110010000: color_data = 108'b111111111111111111111111110111011101111111111111110111011101111111111111110111011101111111111111101010011010;
		12'b101110010001: color_data = 108'b110111011101111111111111100010001001110111011101101010011010111111111111100110011010110111011101100001100110;
		12'b101110010010: color_data = 108'b100010001001110111011101100110011010100110011010100001100110110111011101101110111100101010011010011101111000;
		12'b101110010011: color_data = 108'b100110011010100010001001101010101011101110111100011101111000100110011010110011001101100001100110011101111000;
		12'b101110010100: color_data = 108'b101010101011100110011010101110111100110011001101011101111000101110111100110111011110011101111000100001111001;
		12'b101110010101: color_data = 108'b101110111100101010101011110111011110110111011110100001111001110011001101110111101111011101111000101010001001;
		12'b101110010110: color_data = 108'b110111011110101110111100110111011110110111101111101010001001110111011110111011101111100001111001101010001001;
		12'b101110010111: color_data = 108'b110111011110110111011110111011101110111011101111101010001001110111101111111111111111101010001001110110111100;
		12'b101110011000: color_data = 108'b111011101110110111011110110111011101111111111111110110111100111011101111110111011101101010001001110111011101;
		12'b101110011001: color_data = 108'b110111011101111011101110010101010110110111011101110111011101111111111111011001100111110110111100011001100111;
		12'b101110011010: color_data = 108'b010101010110110111011101010101010110011001100111011001100111110111011101011001101000110111011101010001000101;
		12'b101110011011: color_data = 108'b010101010110010101010110011001100110011001101000010001000101011001100111011101111001011001100111010001000101;
		12'b101110011100: color_data = 108'b011001100110010101010110011001100111011101111001010001000101011001101000011101111001010001000101010101010101;
		12'b101110011101: color_data = 108'b011001100111011001100110011101111000011101111001010101010101011101111001100010001001010001000101011101111000;
		12'b101110011110: color_data = 108'b011101111000011001100111100110011010100010001001011101111000011101111001110011001101010101010101100001100111;
		12'b101110011111: color_data = 108'b100110011010011101111000110011001100110011001101100001100111100010001001111111111111011101111000101010001001;
		12'b101110100000: color_data = 108'b110011001100100110011010111111111111111111111111101010001001110011001101111111111111100001100111111111111111;
		12'b101110100001: color_data = 108'b111111111111110011001100111111111111111111111111111111111111111111111111111111111111101010001001111111111111;
		12'b101110100010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110100011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b101111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111001111: color_data = 108'b111111111111111111111111110111011101111111111111111111111111111111111111111111111111111111111111011101110111;
		12'b101111010000: color_data = 108'b110111011101111111111111101010011010111111111111011101110111111111111111110111011101111111111111010000010001;
		12'b101111010001: color_data = 108'b101010011010110111011101100001100110110111011101010000010001111111111111100010001001011101110111100000000000;
		12'b101111010010: color_data = 108'b100001100110101010011010011101111000100010001001100000000000110111011101100110011010010000010001100001100111;
		12'b101111010011: color_data = 108'b011101111000100001100110011101111000100110011010100001100111100010001001101010101011100000000000011101111000;
		12'b101111010100: color_data = 108'b011101111000011101111000100001111001101010101011011101111000100110011010101110111100100001100111100001100110;
		12'b101111010101: color_data = 108'b100001111001011101111000101010001001101110111100100001100110101010101011110111011110011101111000100100010001;
		12'b101111010110: color_data = 108'b101010001001100001111001101010001001110111011110100100010001101110111100110111011110100001100110100100000001;
		12'b101111010111: color_data = 108'b101010001001101010001001110110111100110111011110100100000001110111011110111011101110100100010001110001110111;
		12'b101111011000: color_data = 108'b110110111100101010001001110111011101111011101110110001110111110111011110110111011101100100000001111011101110;
		12'b101111011001: color_data = 108'b110111011101110110111100011001100111110111011101111011101110111011101110010101010110110001110111100010001001;
		12'b101111011010: color_data = 108'b011001100111110111011101010001000101010101010110100010001001110111011101010101010110111011101110011001010110;
		12'b101111011011: color_data = 108'b010001000101011001100111010001000101010101010110011001010110010101010110011001100110100010001001010101000101;
		12'b101111011100: color_data = 108'b010001000101010001000101010101010101011001100110010101000101010101010110011001100111011001010110010101000101;
		12'b101111011101: color_data = 108'b010101010101010001000101011101111000011001100111010101000101011001100110011101111000010101000101011101111000;
		12'b101111011110: color_data = 108'b011101111000010101010101100001100111011101111000011101111000011001100111100110011010010101000101100000100011;
		12'b101111011111: color_data = 108'b100001100111011101111000101010001001100110011010100000100011011101111000110011001100011101111000101001000100;
		12'b101111100000: color_data = 108'b101010001001100001100111111111111111110011001100101001000100100110011010111111111111100000100011111011101110;
		12'b101111100001: color_data = 108'b111111111111101010001001111111111111111111111111111011101110110011001100111111111111101001000100111011101110;
		12'b101111100010: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111011101110111011101111;
		12'b101111100011: color_data = 108'b111111111111111111111111111111111111111111111111111011101111111111111111111111111111111011101110111111111111;
		12'b101111100100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111111;
		12'b101111100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b101111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110000000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000001111: color_data = 108'b111111111111111111111111011101110111111111111111111111111111111111111111110111011101111111111111011101110111;
		12'b110000010000: color_data = 108'b011101110111111111111111010000010001110111011101011101110111111111111111101010011010111111111111010000010001;
		12'b110000010001: color_data = 108'b010000010001011101110111100000000000101010011010010000010001110111011101100001100110011101110111100000000000;
		12'b110000010010: color_data = 108'b100000000000010000010001100001100111100001100110100000000000101010011010011101111000010000010001100000010001;
		12'b110000010011: color_data = 108'b100001100111100000000000011101111000011101111000100000010001100001100110011101111000100000000000100000010001;
		12'b110000010100: color_data = 108'b011101111000100001100111100001100110011101111000100000010001011101111000100001111001100000010001100100110011;
		12'b110000010101: color_data = 108'b100001100110011101111000100100010001100001111001100100110011011101111000101010001001100000010001101110011010;
		12'b110000010110: color_data = 108'b100100010001100001100110100100000001101010001001101110011010100001111001101010001001100100110011110110111011;
		12'b110000010111: color_data = 108'b100100000001100100010001110001110111101010001001110110111011101010001001110110111100101110011010101110111011;
		12'b110000011000: color_data = 108'b110001110111100100000001111011101110110110111100101110111011101010001001110111011101110110111011100110011010;
		12'b110000011001: color_data = 108'b111011101110110001110111100010001001110111011101100110011010110110111100011001100111101110111011100010001001;
		12'b110000011010: color_data = 108'b100010001001111011101110011001010110011001100111100010001001110111011101010001000101100110011010110000110011;
		12'b110000011011: color_data = 108'b011001010110100010001001010101000101010001000101110000110011011001100111010001000101100010001001100100010001;
		12'b110000011100: color_data = 108'b010101000101011001010110010101000101010001000101100100010001010001000101010101010101110000110011001000100011;
		12'b110000011101: color_data = 108'b010101000101010101000101011101111000010101010101001000100011010001000101011101111000100100010001001100110011;
		12'b110000011110: color_data = 108'b011101111000010101000101100000100011011101111000001100110011010101010101100001100111001000100011010000110100;
		12'b110000011111: color_data = 108'b100000100011011101111000101001000100100001100111010000110100011101111000101010001001001100110011011001010110;
		12'b110000100000: color_data = 108'b101001000100100000100011111011101110101010001001011001010110100001100111111111111111010000110100100110011010;
		12'b110000100001: color_data = 108'b111011101110101001000100111011101110111111111111100110011010101010001001111111111111011001010110100110011010;
		12'b110000100010: color_data = 108'b111011101110111011101110111011101111111111111111100110011010111111111111111111111111100110011010110011001101;
		12'b110000100011: color_data = 108'b111011101111111011101110111111111111111111111111110011001101111111111111111111111111100110011010111111111111;
		12'b110000100100: color_data = 108'b111111111111111011101111111111111111111111111111111111111111111111111111111111111111110011001101111111111111;
		12'b110000100101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000100110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110000101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110001000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110;
		12'b110001001110: color_data = 108'b111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111100110011001;
		12'b110001001111: color_data = 108'b111111111111111111111111011101110111111111111111100110011001111111111111011101110111111011101110011000110011;
		12'b110001010000: color_data = 108'b011101110111111111111111010000010001011101110111011000110011111111111111010000010001100110011001011000000000;
		12'b110001010001: color_data = 108'b010000010001011101110111100000000000010000010001011000000000011101110111100000000000011000110011100000000000;
		12'b110001010010: color_data = 108'b100000000000010000010001100000010001100000000000100000000000010000010001100001100111011000000000100000000000;
		12'b110001010011: color_data = 108'b100000010001100000000000100000010001100001100111100000000000100000000000011101111000100000000000100000010010;
		12'b110001010100: color_data = 108'b100000010001100000010001100100110011011101111000100000010010100001100111100001100110100000000000100101010110;
		12'b110001010101: color_data = 108'b100100110011100000010001101110011010100001100110100101010110011101111000100100010001100000010010101110111100;
		12'b110001010110: color_data = 108'b101110011010100100110011110110111011100100010001101110111100100001100110100100000001100101010110111010001001;
		12'b110001010111: color_data = 108'b110110111011101110011010101110111011100100000001111010001001100100010001110001110111101110111100111001010110;
		12'b110001011000: color_data = 108'b101110111011110110111011100110011010110001110111111001010110100100000001111011101110111010001001101100110100;
		12'b110001011001: color_data = 108'b100110011010101110111011100010001001111011101110101100110100110001110111100010001001111001010110110000110100;
		12'b110001011010: color_data = 108'b100010001001100110011010110000110011100010001001110000110100111011101110011001010110101100110100111000010001;
		12'b110001011011: color_data = 108'b110000110011100010001001100100010001011001010110111000010001100010001001010101000101110000110100110100000000;
		12'b110001011100: color_data = 108'b100100010001110000110011001000100011010101000101110100000000011001010110010101000101111000010001100100010001;
		12'b110001011101: color_data = 108'b001000100011100100010001001100110011010101000101100100010001010101000101011101111000110100000000100100010001;
		12'b110001011110: color_data = 108'b001100110011001000100011010000110100011101111000100100010001010101000101100000100011100100010001010100100010;
		12'b110001011111: color_data = 108'b010000110100001100110011011001010110100000100011010100100010011101111000101001000100100100010001001101000100;
		12'b110001100000: color_data = 108'b011001010110010000110100100110011010101001000100001101000100100000100011111011101110010100100010010001010101;
		12'b110001100001: color_data = 108'b100110011010011001010110100110011010111011101110010001010101101001000100111011101110001101000100010001010101;
		12'b110001100010: color_data = 108'b100110011010100110011010110011001101111011101110010001010101111011101110111011101111010001010101100001100110;
		12'b110001100011: color_data = 108'b110011001101100110011010111111111111111011101111100001100110111011101110111111111111010001010101110001110111;
		12'b110001100100: color_data = 108'b111111111111110011001101111111111111111111111111110001110111111011101111111111111111100001100110110001110111;
		12'b110001100101: color_data = 108'b111111111111111111111111111111111111111111111111110001110111111111111111111111111111110001110111111011011101;
		12'b110001100110: color_data = 108'b111111111111111111111111111111111111111111111111111011011101111111111111111111111111110001110111111111111111;
		12'b110001100111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011101111111111111;
		12'b110001101000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001101001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110001101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110010000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010001101: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111111111111111111111111111110111011101;
		12'b110010001110: color_data = 108'b111011101110111111111111100110011001111111111111110111011101111111111111111111111111111111111111001100110011;
		12'b110010001111: color_data = 108'b100110011001111011101110011000110011111111111111001100110011111111111111011101110111110111011101011000000000;
		12'b110010010000: color_data = 108'b011000110011100110011001011000000000011101110111011000000000111111111111010000010001001100110011100100000000;
		12'b110010010001: color_data = 108'b011000000000011000110011100000000000010000010001100100000000011101110111100000000000011000000000100000000000;
		12'b110010010010: color_data = 108'b100000000000011000000000100000000000100000000000100000000000010000010001100000010001100100000000100000000000;
		12'b110010010011: color_data = 108'b100000000000100000000000100000010010100000010001100000000000100000000000100000010001100000000000100001000100;
		12'b110010010100: color_data = 108'b100000010010100000000000100101010110100000010001100001000100100000010001100100110011100000000000100110001001;
		12'b110010010101: color_data = 108'b100101010110100000010010101110111100100100110011100110001001100000010001101110011010100001000100110010001001;
		12'b110010010110: color_data = 108'b101110111100100101010110111010001001101110011010110010001001100100110011110110111011100110001001111100100010;
		12'b110010010111: color_data = 108'b111010001001101110111100111001010110110110111011111100100010101110011010101110111011110010001001111100000000;
		12'b110010011000: color_data = 108'b111001010110111010001001101100110100101110111011111100000000110110111011100110011010111100100010111100000000;
		12'b110010011001: color_data = 108'b101100110100111001010110110000110100100110011010111100000000101110111011100010001001111100000000111100000000;
		12'b110010011010: color_data = 108'b110000110100101100110100111000010001100010001001111100000000100110011010110000110011111100000000111100000000;
		12'b110010011011: color_data = 108'b111000010001110000110100110100000000110000110011111100000000100010001001100100010001111100000000111100000000;
		12'b110010011100: color_data = 108'b110100000000111000010001100100010001100100010001111100000000110000110011001000100011111100000000111100000000;
		12'b110010011101: color_data = 108'b100100010001110100000000100100010001001000100011111100000000100100010001001100110011111100000000111100000000;
		12'b110010011110: color_data = 108'b100100010001100100010001010100100010001100110011111100000000001000100011010000110100111100000000100100010001;
		12'b110010011111: color_data = 108'b010100100010100100010001001101000100010000110100100100010001001100110011011001010110111100000000010100010001;
		12'b110010100000: color_data = 108'b001101000100010100100010010001010101011001010110010100010001010000110100100110011010100100010001010100010001;
		12'b110010100001: color_data = 108'b010001010101001101000100010001010101100110011010010100010001011001010110100110011010010100010001010100010001;
		12'b110010100010: color_data = 108'b010001010101010001010101100001100110100110011010010100010001100110011010110011001101010100010001011000000000;
		12'b110010100011: color_data = 108'b100001100110010001010101110001110111110011001101011000000000100110011010111111111111010100010001011100000000;
		12'b110010100100: color_data = 108'b110001110111100001100110110001110111111111111111011100000000110011001101111111111111011000000000011100000000;
		12'b110010100101: color_data = 108'b110001110111110001110111111011011101111111111111011100000000111111111111111111111111011100000000110010011001;
		12'b110010100110: color_data = 108'b111011011101110001110111111111111111111111111111110010011001111111111111111111111111011100000000111011001100;
		12'b110010100111: color_data = 108'b111111111111111011011101111111111111111111111111111011001100111111111111111111111111110010011001111011001100;
		12'b110010101000: color_data = 108'b111111111111111111111111111111111111111111111111111011001100111111111111111111111111111011001100111111101110;
		12'b110010101001: color_data = 108'b111111111111111111111111111111111111111111111111111111101110111111111111111111111111111011001100111111111111;
		12'b110010101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111111;
		12'b110010101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110010101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110011000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011001101: color_data = 108'b111111111111111111111111110111011101111111111111111111111111111111111111111011101110111111111111110111011101;
		12'b110011001110: color_data = 108'b110111011101111111111111001100110011111011101110110111011101111111111111100110011001111111111111001100110011;
		12'b110011001111: color_data = 108'b001100110011110111011101011000000000100110011001001100110011111011101110011000110011110111011101011000000000;
		12'b110011010000: color_data = 108'b011000000000001100110011100100000000011000110011011000000000100110011001011000000000001100110011100000000000;
		12'b110011010001: color_data = 108'b100100000000011000000000100000000000011000000000100000000000011000110011100000000000011000000000100000000000;
		12'b110011010010: color_data = 108'b100000000000100100000000100000000000100000000000100000000000011000000000100000000000100000000000100000000000;
		12'b110011010011: color_data = 108'b100000000000100000000000100001000100100000000000100000000000100000000000100000010010100000000000100001000100;
		12'b110011010100: color_data = 108'b100001000100100000000000100110001001100000010010100001000100100000000000100101010110100000000000100101100111;
		12'b110011010101: color_data = 108'b100110001001100001000100110010001001100101010110100101100111100000010010101110111100100001000100111100000001;
		12'b110011010110: color_data = 108'b110010001001100110001001111100100010101110111100111100000001100101010110111010001001100101100111111100000000;
		12'b110011010111: color_data = 108'b111100100010110010001001111100000000111010001001111100000000101110111100111001010110111100000001111100000000;
		12'b110011011000: color_data = 108'b111100000000111100100010111100000000111001010110111100000000111010001001101100110100111100000000111100000000;
		12'b110011011001: color_data = 108'b111100000000111100000000111100000000101100110100111100000000111001010110110000110100111100000000111100000000;
		12'b110011011010: color_data = 108'b111100000000111100000000111100000000110000110100111100000000101100110100111000010001111100000000111100000000;
		12'b110011011011: color_data = 108'b111100000000111100000000111100000000111000010001111100000000110000110100110100000000111100000000111100000000;
		12'b110011011100: color_data = 108'b111100000000111100000000111100000000110100000000111100000000111000010001100100010001111100000000111100000000;
		12'b110011011101: color_data = 108'b111100000000111100000000111100000000100100010001111100000000110100000000100100010001111100000000111100000000;
		12'b110011011110: color_data = 108'b111100000000111100000000100100010001100100010001111100000000100100010001010100100010111100000000111100000000;
		12'b110011011111: color_data = 108'b100100010001111100000000010100010001010100100010111100000000100100010001001101000100111100000000111000000000;
		12'b110011100000: color_data = 108'b010100010001100100010001010100010001001101000100111000000000010100100010010001010101111100000000111000000000;
		12'b110011100001: color_data = 108'b010100010001010100010001010100010001010001010101111000000000001101000100010001010101111000000000111000000000;
		12'b110011100010: color_data = 108'b010100010001010100010001011000000000010001010101111000000000010001010101100001100110111000000000100000010001;
		12'b110011100011: color_data = 108'b011000000000010100010001011100000000100001100110100000010001010001010101110001110111111000000000001000100010;
		12'b110011100100: color_data = 108'b011100000000011000000000011100000000110001110111001000100010100001100110110001110111100000010001001000100010;
		12'b110011100101: color_data = 108'b011100000000011100000000110010011001110001110111001000100010110001110111111011011101001000100010011100010001;
		12'b110011100110: color_data = 108'b110010011001011100000000111011001100111011011101011100010001110001110111111111111111001000100010100100000000;
		12'b110011100111: color_data = 108'b111011001100110010011001111011001100111111111111100100000000111011011101111111111111011100010001101000110011;
		12'b110011101000: color_data = 108'b111011001100111011001100111111101110111111111111101000110011111111111111111111111111100100000000111011101110;
		12'b110011101001: color_data = 108'b111111101110111011001100111111111111111111111111111011101110111111111111111111111111101000110011111111111111;
		12'b110011101010: color_data = 108'b111111111111111111101110111111111111111111111111111111111111111111111111111111111111111011101110111111111111;
		12'b110011101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110011101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110100000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100001101: color_data = 108'b111111111111111111111111110111011101111111111111111111111111111111111111110111011101111111111111110111011101;
		12'b110100001110: color_data = 108'b110111011101111111111111001100110011110111011101110111011101111111111111001100110011111111111111001100110011;
		12'b110100001111: color_data = 108'b001100110011110111011101011000000000001100110011001100110011110111011101011000000000110111011101001100010001;
		12'b110100010000: color_data = 108'b011000000000001100110011100000000000011000000000001100010001001100110011100100000000001100110011001100010001;
		12'b110100010001: color_data = 108'b100000000000011000000000100000000000100100000000001100010001011000000000100000000000001100010001001100010001;
		12'b110100010010: color_data = 108'b100000000000100000000000100000000000100000000000001100010001100100000000100000000000001100010001001100010001;
		12'b110100010011: color_data = 108'b100000000000100000000000100001000100100000000000001100010001100000000000100001000100001100010001001100100010;
		12'b110100010100: color_data = 108'b100001000100100000000000100101100111100001000100001100100010100000000000100110001001001100010001010000110011;
		12'b110100010101: color_data = 108'b100101100111100001000100111100000001100110001001010000110011100001000100110010001001001100100010010100010001;
		12'b110100010110: color_data = 108'b111100000001100101100111111100000000110010001001010100010001100110001001111100100010010000110011010100010001;
		12'b110100010111: color_data = 108'b111100000000111100000001111100000000111100100010010100010001110010001001111100000000010100010001010100010001;
		12'b110100011000: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100100010111100000000010100010001010100010001;
		12'b110100011001: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100000000111100000000010100010001010100010001;
		12'b110100011010: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100000000111100000000010100010001010100010001;
		12'b110100011011: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100000000111100000000010100010001010100010001;
		12'b110100011100: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100000000111100000000010100010001010100010001;
		12'b110100011101: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100000000111100000000010100010001010100010001;
		12'b110100011110: color_data = 108'b111100000000111100000000111100000000111100000000010100010001111100000000100100010001010100010001010100010001;
		12'b110100011111: color_data = 108'b111100000000111100000000111000000000100100010001010100010001111100000000010100010001010100010001010100010001;
		12'b110100100000: color_data = 108'b111000000000111100000000111000000000010100010001010100010001100100010001010100010001010100010001010100010001;
		12'b110100100001: color_data = 108'b111000000000111000000000111000000000010100010001010100010001010100010001010100010001010100010001010100010001;
		12'b110100100010: color_data = 108'b111000000000111000000000100000010001010100010001010100010001010100010001011000000000010100010001001100010001;
		12'b110100100011: color_data = 108'b100000010001111000000000001000100010011000000000001100010001010100010001011100000000010100010001001000100010;
		12'b110100100100: color_data = 108'b001000100010100000010001001000100010011100000000001000100010011000000000011100000000001100010001001000100010;
		12'b110100100101: color_data = 108'b001000100010001000100010011100010001011100000000001000100010011100000000110010011001001000100010001100010001;
		12'b110100100110: color_data = 108'b011100010001001000100010100100000000110010011001001100010001011100000000111011001100001000100010001100010001;
		12'b110100100111: color_data = 108'b100100000000011100010001101000110011111011001100001100010001110010011001111011001100001100010001010100110011;
		12'b110100101000: color_data = 108'b101000110011100100000000111011101110111011001100010100110011111011001100111111101110001100010001111011101110;
		12'b110100101001: color_data = 108'b111011101110101000110011111111111111111111101110111011101110111011001100111111111111010100110011111111111111;
		12'b110100101010: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111111101110111111111111111011101110111111111111;
		12'b110100101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110100101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110101000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101001101: color_data = 108'b111111111111111111111111110111011101111111111111111111111111111111111111110111011101111111111111111011101110;
		12'b110101001110: color_data = 108'b110111011101111111111111001100110011110111011101111011101110111111111111001100110011111111111111100010001000;
		12'b110101001111: color_data = 108'b001100110011110111011101001100010001001100110011100010001000110111011101011000000000111011101110011101110111;
		12'b110101010000: color_data = 108'b001100010001001100110011001100010001011000000000011101110111001100110011100000000000100010001000011101110111;
		12'b110101010001: color_data = 108'b001100010001001100010001001100010001100000000000011101110111011000000000100000000000011101110111011101110111;
		12'b110101010010: color_data = 108'b001100010001001100010001001100010001100000000000011101110111100000000000100000000000011101110111011101110111;
		12'b110101010011: color_data = 108'b001100010001001100010001001100100010100000000000011101110111100000000000100001000100011101110111011101110111;
		12'b110101010100: color_data = 108'b001100100010001100010001010000110011100001000100011101110111100000000000100101100111011101110111011101110111;
		12'b110101010101: color_data = 108'b010000110011001100100010010100010001100101100111011101110111100001000100111100000001011101110111011101110111;
		12'b110101010110: color_data = 108'b010100010001010000110011010100010001111100000001011101110111100101100111111100000000011101110111011101110111;
		12'b110101010111: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000001111100000000011101110111011101110111;
		12'b110101011000: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011001: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011010: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011011: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011100: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011101: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011110: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111100000000011101110111011101110111;
		12'b110101011111: color_data = 108'b010100010001010100010001010100010001111100000000011101110111111100000000111000000000011101110111011101110111;
		12'b110101100000: color_data = 108'b010100010001010100010001010100010001111000000000011101110111111100000000111000000000011101110111011101110111;
		12'b110101100001: color_data = 108'b010100010001010100010001010100010001111000000000011101110111111000000000111000000000011101110111011101110111;
		12'b110101100010: color_data = 108'b010100010001010100010001001100010001111000000000011101110111111000000000100000010001011101110111011101110111;
		12'b110101100011: color_data = 108'b001100010001010100010001001000100010100000010001011101110111111000000000001000100010011101110111011101110111;
		12'b110101100100: color_data = 108'b001000100010001100010001001000100010001000100010011101110111100000010001001000100010011101110111011101110111;
		12'b110101100101: color_data = 108'b001000100010001000100010001100010001001000100010011101110111001000100010011100010001011101110111011101110111;
		12'b110101100110: color_data = 108'b001100010001001000100010001100010001011100010001011101110111001000100010100100000000011101110111011101110111;
		12'b110101100111: color_data = 108'b001100010001001100010001010100110011100100000000011101110111011100010001101000110011011101110111100110011001;
		12'b110101101000: color_data = 108'b010100110011001100010001111011101110101000110011100110011001100100000000111011101110011101110111111011101110;
		12'b110101101001: color_data = 108'b111011101110010100110011111111111111111011101110111011101110101000110011111111111111100110011001111111111111;
		12'b110101101010: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111011101110111111111111111011101110111111111111;
		12'b110101101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110101101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110110000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110001101: color_data = 108'b111111111111111111111111111011101110111111111111111111111111111111111111110111011101111111111111111111111111;
		12'b110110001110: color_data = 108'b111011101110111111111111100010001000110111011101111111111111111111111111001100110011111111111111111111111111;
		12'b110110001111: color_data = 108'b100010001000111011101110011101110111001100110011111111111111110111011101001100010001111111111111111111111111;
		12'b110110010000: color_data = 108'b011101110111100010001000011101110111001100010001111111111111001100110011001100010001111111111111111111111111;
		12'b110110010001: color_data = 108'b011101110111011101110111011101110111001100010001111111111111001100010001001100010001111111111111111111111111;
		12'b110110010010: color_data = 108'b011101110111011101110111011101110111001100010001111111111111001100010001001100010001111111111111111111111111;
		12'b110110010011: color_data = 108'b011101110111011101110111011101110111001100010001111111111111001100010001001100100010111111111111111111111111;
		12'b110110010100: color_data = 108'b011101110111011101110111011101110111001100100010111111111111001100010001010000110011111111111111111111111111;
		12'b110110010101: color_data = 108'b011101110111011101110111011101110111010000110011111111111111001100100010010100010001111111111111111111111111;
		12'b110110010110: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010000110011010100010001111111111111111111111111;
		12'b110110010111: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011000: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011001: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011010: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011011: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011100: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011101: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011110: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110011111: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110100000: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110100001: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001010100010001111111111111111111111111;
		12'b110110100010: color_data = 108'b011101110111011101110111011101110111010100010001111111111111010100010001001100010001111111111111111111111111;
		12'b110110100011: color_data = 108'b011101110111011101110111011101110111001100010001111111111111010100010001001000100010111111111111111111111111;
		12'b110110100100: color_data = 108'b011101110111011101110111011101110111001000100010111111111111001100010001001000100010111111111111111111111111;
		12'b110110100101: color_data = 108'b011101110111011101110111011101110111001000100010111111111111001000100010001100010001111111111111111111111111;
		12'b110110100110: color_data = 108'b011101110111011101110111011101110111001100010001111111111111001000100010001100010001111111111111111111111111;
		12'b110110100111: color_data = 108'b011101110111011101110111100110011001001100010001111111111111001100010001010100110011111111111111111111111111;
		12'b110110101000: color_data = 108'b100110011001011101110111111011101110010100110011111111111111001100010001111011101110111111111111111111111111;
		12'b110110101001: color_data = 108'b111011101110100110011001111111111111111011101110111111111111010100110011111111111111111111111111111111111111;
		12'b110110101010: color_data = 108'b111111111111111011101110111111111111111111111111111111111111111011101110111111111111111111111111111111111111;
		12'b110110101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110110101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		12'b110111000000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000110: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111000111: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111001000: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111001001: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111001010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111001011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111001100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111001101: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111;
		12'b110111001110: color_data = 108'b111111111111111111111111111111111111111011101110111111111111111111111111100010001000111111111111111111111111;
		12'b110111001111: color_data = 108'b111111111111111111111111111111111111100010001000111111111111111011101110011101110111111111111111111111111111;
		12'b110111010000: color_data = 108'b111111111111111111111111111111111111011101110111111111111111100010001000011101110111111111111111111111111111;
		12'b110111010001: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111010010: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111010011: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111010100: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111010101: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111010110: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111010111: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011000: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011001: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011010: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011011: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011100: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011101: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011110: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111011111: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100000: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100001: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100010: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100011: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100100: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100101: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100110: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111011101110111111111111111111111111111;
		12'b110111100111: color_data = 108'b111111111111111111111111111111111111011101110111111111111111011101110111100110011001111111111111111111111111;
		12'b110111101000: color_data = 108'b111111111111111111111111111111111111100110011001111111111111011101110111111011101110111111111111111111111111;
		12'b110111101001: color_data = 108'b111111111111111111111111111111111111111011101110111111111111100110011001111111111111111111111111111111111111;
		12'b110111101010: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111011101110111111111111111111111111111111111111;
		12'b110111101011: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		12'b110111101100: color_data = 108'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

		default: color_data = 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase
endmodule